/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
Control_Alu
**
**
**
*****************************************************************************/
module
Control_Alu(
Opcode,
aluop,
funct
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[5:0]
Opcode;
input
[5:0]
funct;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
[3:0]
aluop;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[3:0]
s_logisimBus10;
wire
[3:0]
s_logisimBus11;
wire
[3:0]
s_logisimBus12;
wire
[5:0]
s_logisimBus13;
wire
[3:0]
s_logisimBus19;
wire
[5:0]
s_logisimBus20;
wire
[3:0]
s_logisimBus24;
wire
[3:0]
s_logisimBus25;
wire
[3:0]
s_logisimBus26;
wire
[3:0]
s_logisimBus27;
wire
[3:0]
s_logisimBus30;
wire
[5:0]
s_logisimBus32;
wire
[5:0]
s_logisimBus33;
wire
[5:0]
s_logisimBus34;
wire
[3:0]
s_logisimBus37;
wire
[3:0]
s_logisimBus38;
wire
[5:0]
s_logisimBus4;
wire
[3:0]
s_logisimBus43;
wire
[5:0]
s_logisimBus45;
wire
[5:0]
s_logisimBus47;
wire
[3:0]
s_logisimBus48;
wire
s_logisimNet0;
wire
s_logisimNet1;
wire
s_logisimNet14;
wire
s_logisimNet15;
wire
s_logisimNet16;
wire
s_logisimNet17;
wire
s_logisimNet18;
wire
s_logisimNet2;
wire
s_logisimNet21;
wire
s_logisimNet22;
wire
s_logisimNet23;
wire
s_logisimNet28;
wire
s_logisimNet29;
wire
s_logisimNet3;
wire
s_logisimNet31;
wire
s_logisimNet35;
wire
s_logisimNet36;
wire
s_logisimNet39;
wire
s_logisimNet40;
wire
s_logisimNet41;
wire
s_logisimNet42;
wire
s_logisimNet44;
wire
s_logisimNet46;
wire
s_logisimNet49;
wire
s_logisimNet5;
wire
s_logisimNet6;
wire
s_logisimNet7;
wire
s_logisimNet8;
wire
s_logisimNet9;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus13[5:0]
=
Opcode;
assign
s_logisimBus4[5:0]
=
funct;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
aluop
=
s_logisimBus38[3:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus47[5:0]
=
{2'b00,
4'h2};
assign
s_logisimBus37[3:0]
=
4'h2;
assign
s_logisimBus32[5:0]
=
{2'b01,
4'hA};
assign
s_logisimBus25[3:0]
=
4'h3;
assign
s_logisimBus20[5:0]
=
{2'b00,
4'h0};
assign
s_logisimBus27[3:0]
=
4'h1;
assign
s_logisimBus43[3:0]
=
4'h0;
assign
s_logisimBus48[3:0]
=
4'h9;
assign
s_logisimBus19[3:0]
=
4'h0;
assign
s_logisimBus34[5:0]
=
{2'b00,
4'h8};
assign
s_logisimBus45[5:0]
=
{2'b00,
4'h0};
assign
s_logisimBus33[5:0]
=
{2'b01,
4'hC};
assign
s_logisimNet9
=
~s_logisimNet15;
assign
s_logisimNet22
=
~s_logisimBus4[5];
assign
s_logisimNet41
=
~s_logisimBus4[5];
assign
s_logisimNet23
=
~s_logisimBus4[1];
assign
s_logisimNet36
=
~s_logisimBus4[0];
assign
s_logisimNet6
=
~s_logisimBus4[1];
assign
s_logisimNet7
=
~s_logisimBus4[2];
assign
s_logisimNet42
=
~s_logisimBus4[0];
assign
s_logisimNet16
=
~s_logisimNet46;
assign
s_logisimBus30[3]
=
~s_logisimBus4[5];
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
AND_GATE
#(.BubblesMask(2'b00))
GATES_1
(.input1(s_logisimBus4[1]),
.input2(s_logisimBus4[2]),
.result(s_logisimBus30[1]));
AND_GATE
#(.BubblesMask(2'b00))
GATES_2
(.input1(s_logisimBus4[2]),
.input2(s_logisimBus4[5]),
.result(s_logisimBus30[2]));
AND_GATE
#(.BubblesMask(2'b00))
GATES_3
(.input1(s_logisimNet9),
.input2(s_logisimNet16),
.result(s_logisimNet35));
AND_GATE_4_INPUTS
#(.BubblesMask(4'h0))
GATES_4
(.input1(s_logisimBus4[2]),
.input2(s_logisimNet22),
.input3(s_logisimBus4[1]),
.input4(s_logisimBus4[0]),
.result(s_logisimNet17));
AND_GATE_4_INPUTS
#(.BubblesMask(4'h0))
GATES_5
(.input1(s_logisimBus4[2]),
.input2(s_logisimNet41),
.input3(s_logisimNet23),
.input4(s_logisimNet36),
.result(s_logisimNet40));
AND_GATE_4_INPUTS
#(.BubblesMask(4'h0))
GATES_6
(.input1(s_logisimBus4[2]),
.input2(s_logisimBus4[5]),
.input3(s_logisimNet6),
.input4(s_logisimBus4[0]),
.result(s_logisimNet29));
AND_GATE_4_INPUTS
#(.BubblesMask(4'h0))
GATES_7
(.input1(s_logisimBus4[5]),
.input2(s_logisimNet7),
.input3(s_logisimBus4[1]),
.input4(s_logisimNet42),
.result(s_logisimNet18));
OR_GATE_4_INPUTS
#(.BubblesMask(4'h0))
GATES_8
(.input1(s_logisimNet17),
.input2(s_logisimNet40),
.input3(s_logisimNet29),
.input4(s_logisimNet18),
.result(s_logisimBus30[0]));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_9
(.enable(1'b1),
.muxIn_0(s_logisimBus30[3:0]),
.muxIn_1(s_logisimBus37[3:0]),
.muxOut(s_logisimBus10[3:0]),
.sel(s_logisimNet44));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_10
(.enable(1'b1),
.muxIn_0(s_logisimBus10[3:0]),
.muxIn_1(s_logisimBus25[3:0]),
.muxOut(s_logisimBus26[3:0]),
.sel(s_logisimNet39));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_11
(.enable(1'b1),
.muxIn_0(s_logisimBus26[3:0]),
.muxIn_1(s_logisimBus48[3:0]),
.muxOut(s_logisimBus24[3:0]),
.sel(s_logisimNet14));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_12
(.enable(1'b1),
.muxIn_0(s_logisimBus27[3:0]),
.muxIn_1(s_logisimBus43[3:0]),
.muxOut(s_logisimBus11[3:0]),
.sel(s_logisimBus13[5]));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_13
(.enable(1'b1),
.muxIn_0(s_logisimBus24[3:0]),
.muxIn_1(s_logisimBus12[3:0]),
.muxOut(s_logisimBus38[3:0]),
.sel(s_logisimNet35));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_14
(.enable(1'b1),
.muxIn_0(s_logisimBus11[3:0]),
.muxIn_1(s_logisimBus19[3:0]),
.muxOut(s_logisimBus12[3:0]),
.sel(s_logisimNet3));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_15
(.aEqualsB(s_logisimNet44),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus4[5:0]),
.dataB(s_logisimBus47[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_16
(.aEqualsB(s_logisimNet39),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus32[5:0]),
.dataB(s_logisimBus4[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_17
(.aEqualsB(s_logisimNet14),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus20[5:0]),
.dataB(s_logisimBus4[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_18
(.aEqualsB(s_logisimNet3),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus34[5:0]),
.dataB(s_logisimBus13[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_19
(.aEqualsB(s_logisimNet15),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus13[5:0]),
.dataB(s_logisimBus45[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_20
(.aEqualsB(s_logisimNet46),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus13[5:0]),
.dataB(s_logisimBus33[5:0]));
endmodule