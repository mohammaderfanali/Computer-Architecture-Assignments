/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
AND_GATE_4_INPUTS
**
**
**
*****************************************************************************/
module
AND_GATE_4_INPUTS(
input1,
input2,
input3,
input4,
result
);
/*******************************************************************************
**
Here
all
module
parameters
are
defined
with
a
dummy
value
**
*******************************************************************************/
parameter
[64:0]
BubblesMask
=
1;
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
input1;
input
input2;
input
input3;
input
input4;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
result;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
s_realInput1;
wire
s_realInput2;
wire
s_realInput3;
wire
s_realInput4;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
the
bubbles
are
processed
**
*******************************************************************************/
assign
s_realInput1
=
(BubblesMask[0]
==
1'b0)
?
input1
:
~input1;
assign
s_realInput2
=
(BubblesMask[1]
==
1'b0)
?
input2
:
~input2;
assign
s_realInput3
=
(BubblesMask[2]
==
1'b0)
?
input3
:
~input3;
assign
s_realInput4
=
(BubblesMask[3]
==
1'b0)
?
input4
:
~input4;
/*******************************************************************************
**
Here
the
functionality
is
defined
**
*******************************************************************************/
assign
result
=
s_realInput1&
s_realInput2&
s_realInput3&
s_realInput4;
endmodule