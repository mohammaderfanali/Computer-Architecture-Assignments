/******************************************************************************
 ** Logisim-evolution goes FPGA automatic generated Verilog code             **
 ** https://github.com/logisim-evolution/                                    **
 **                                                                          **
 ** Component : regfile                                                      **
 **                                                                          **
 *****************************************************************************/

module regfile( Aread0,
                Aread1,
                Awrite,
                Dread0,
                Dread1,
                Dwrite,
                R1,
                R10,
                R11,
                R12,
                R13,
                R14,
                R15,
                R16,
                R17,
                R18,
                R19,
                R2,
                R20,
                R21,
                R22,
                R23,
                R24,
                R25,
                R26,
                R27,
                R28,
                R29,
                R3,
                R30,
                R31,
                R4,
                R5,
                R6,
                R7,
                R8,
                R9,
                clk,
                rst );

   /*******************************************************************************
   ** The inputs are defined here                                                **
   *******************************************************************************/
   input [4:0]  Aread0;
   input [4:0]  Aread1;
   input [4:0]  Awrite;
   input [31:0] Dwrite;
   input        clk;
   input        rst;

   /*******************************************************************************
   ** The outputs are defined here                                               **
   *******************************************************************************/
   output [31:0] Dread0;
   output [31:0] Dread1;
   output [31:0] R1;
   output [31:0] R10;
   output [31:0] R11;
   output [31:0] R12;
   output [31:0] R13;
   output [31:0] R14;
   output [31:0] R15;
   output [31:0] R16;
   output [31:0] R17;
   output [31:0] R18;
   output [31:0] R19;
   output [31:0] R2;
   output [31:0] R20;
   output [31:0] R21;
   output [31:0] R22;
   output [31:0] R23;
   output [31:0] R24;
   output [31:0] R25;
   output [31:0] R26;
   output [31:0] R27;
   output [31:0] R28;
   output [31:0] R29;
   output [31:0] R3;
   output [31:0] R30;
   output [31:0] R31;
   output [31:0] R4;
   output [31:0] R5;
   output [31:0] R6;
   output [31:0] R7;
   output [31:0] R8;
   output [31:0] R9;

   /*******************************************************************************
   ** The wires are defined here                                                 **
   *******************************************************************************/
   wire [31:0] s_logisimBus0;
   wire [31:0] s_logisimBus1;
   wire [31:0] s_logisimBus10;
   wire [31:0] s_logisimBus12;
   wire [31:0] s_logisimBus14;
   wire [4:0]  s_logisimBus17;
   wire [31:0] s_logisimBus19;
   wire [31:0] s_logisimBus2;
   wire [31:0] s_logisimBus22;
   wire [31:0] s_logisimBus23;
   wire [31:0] s_logisimBus24;
   wire [31:0] s_logisimBus27;
   wire [31:0] s_logisimBus28;
   wire [31:0] s_logisimBus29;
   wire [31:0] s_logisimBus31;
   wire [31:0] s_logisimBus32;
   wire [31:0] s_logisimBus33;
   wire [31:0] s_logisimBus35;
   wire [31:0] s_logisimBus36;
   wire [4:0]  s_logisimBus37;
   wire [31:0] s_logisimBus38;
   wire [31:0] s_logisimBus39;
   wire [31:0] s_logisimBus40;
   wire [31:0] s_logisimBus41;
   wire [31:0] s_logisimBus42;
   wire [31:0] s_logisimBus43;
   wire [31:0] s_logisimBus44;
   wire [31:0] s_logisimBus45;
   wire [31:0] s_logisimBus46;
   wire [31:0] s_logisimBus47;
   wire [31:0] s_logisimBus49;
   wire [31:0] s_logisimBus50;
   wire [31:0] s_logisimBus52;
   wire [31:0] s_logisimBus53;
   wire [31:0] s_logisimBus54;
   wire [4:0]  s_logisimBus55;
   wire [31:0] s_logisimBus56;
   wire [31:0] s_logisimBus58;
   wire [31:0] s_logisimBus59;
   wire [31:0] s_logisimBus61;
   wire [31:0] s_logisimBus62;
   wire [31:0] s_logisimBus63;
   wire [31:0] s_logisimBus67;
   wire [31:0] s_logisimBus68;
   wire [31:0] s_logisimBus7;
   wire [31:0] s_logisimBus70;
   wire [31:0] s_logisimBus71;
   wire [31:0] s_logisimBus72;
   wire [31:0] s_logisimBus73;
   wire [31:0] s_logisimBus8;
   wire        s_logisimNet100;
   wire        s_logisimNet101;
   wire        s_logisimNet102;
   wire        s_logisimNet103;
   wire        s_logisimNet104;
   wire        s_logisimNet105;
   wire        s_logisimNet106;
   wire        s_logisimNet107;
   wire        s_logisimNet108;
   wire        s_logisimNet109;
   wire        s_logisimNet11;
   wire        s_logisimNet110;
   wire        s_logisimNet111;
   wire        s_logisimNet112;
   wire        s_logisimNet113;
   wire        s_logisimNet114;
   wire        s_logisimNet115;
   wire        s_logisimNet116;
   wire        s_logisimNet117;
   wire        s_logisimNet118;
   wire        s_logisimNet119;
   wire        s_logisimNet120;
   wire        s_logisimNet121;
   wire        s_logisimNet122;
   wire        s_logisimNet123;
   wire        s_logisimNet124;
   wire        s_logisimNet125;
   wire        s_logisimNet126;
   wire        s_logisimNet127;
   wire        s_logisimNet128;
   wire        s_logisimNet129;
   wire        s_logisimNet13;
   wire        s_logisimNet130;
   wire        s_logisimNet131;
   wire        s_logisimNet132;
   wire        s_logisimNet133;
   wire        s_logisimNet134;
   wire        s_logisimNet135;
   wire        s_logisimNet136;
   wire        s_logisimNet137;
   wire        s_logisimNet15;
   wire        s_logisimNet16;
   wire        s_logisimNet18;
   wire        s_logisimNet20;
   wire        s_logisimNet21;
   wire        s_logisimNet25;
   wire        s_logisimNet26;
   wire        s_logisimNet3;
   wire        s_logisimNet30;
   wire        s_logisimNet34;
   wire        s_logisimNet5;
   wire        s_logisimNet51;
   wire        s_logisimNet6;
   wire        s_logisimNet64;
   wire        s_logisimNet66;
   wire        s_logisimNet74;
   wire        s_logisimNet75;
   wire        s_logisimNet76;
   wire        s_logisimNet77;
   wire        s_logisimNet78;
   wire        s_logisimNet79;
   wire        s_logisimNet80;
   wire        s_logisimNet81;
   wire        s_logisimNet82;
   wire        s_logisimNet83;
   wire        s_logisimNet84;
   wire        s_logisimNet85;
   wire        s_logisimNet86;
   wire        s_logisimNet87;
   wire        s_logisimNet88;
   wire        s_logisimNet89;
   wire        s_logisimNet9;
   wire        s_logisimNet90;
   wire        s_logisimNet91;
   wire        s_logisimNet92;
   wire        s_logisimNet93;
   wire        s_logisimNet94;
   wire        s_logisimNet95;
   wire        s_logisimNet96;
   wire        s_logisimNet97;
   wire        s_logisimNet98;
   wire        s_logisimNet99;

   /*******************************************************************************
   ** The module functionality is described here                                 **
   *******************************************************************************/

   /*******************************************************************************
   ** Here all input connections are defined                                     **
   *******************************************************************************/
   assign s_logisimBus17[4:0]  = Awrite;
   assign s_logisimBus37[4:0]  = Aread0;
   assign s_logisimBus55[4:0]  = Aread1;
   assign s_logisimBus73[31:0] = Dwrite;
   assign s_logisimNet3        = clk;
   assign s_logisimNet6        = rst;

   /*******************************************************************************
   ** Here all output connections are defined                                    **
   *******************************************************************************/
   assign Dread0 = s_logisimBus70[31:0];
   assign Dread1 = s_logisimBus63[31:0];
   assign R1     = s_logisimBus43[31:0];
   assign R10    = s_logisimBus44[31:0];
   assign R11    = s_logisimBus54[31:0];
   assign R12    = s_logisimBus14[31:0];
   assign R13    = s_logisimBus24[31:0];
   assign R14    = s_logisimBus45[31:0];
   assign R15    = s_logisimBus56[31:0];
   assign R16    = s_logisimBus2[31:0];
   assign R17    = s_logisimBus32[31:0];
   assign R18    = s_logisimBus1[31:0];
   assign R19    = s_logisimBus31[31:0];
   assign R2     = s_logisimBus27[31:0];
   assign R20    = s_logisimBus19[31:0];
   assign R21    = s_logisimBus42[31:0];
   assign R22    = s_logisimBus53[31:0];
   assign R23    = s_logisimBus62[31:0];
   assign R24    = s_logisimBus7[31:0];
   assign R25    = s_logisimBus33[31:0];
   assign R26    = s_logisimBus49[31:0];
   assign R27    = s_logisimBus28[31:0];
   assign R28    = s_logisimBus29[31:0];
   assign R29    = s_logisimBus35[31:0];
   assign R3     = s_logisimBus46[31:0];
   assign R30    = s_logisimBus50[31:0];
   assign R31    = s_logisimBus59[31:0];
   assign R4     = s_logisimBus58[31:0];
   assign R5     = s_logisimBus12[31:0];
   assign R6     = s_logisimBus40[31:0];
   assign R7     = s_logisimBus23[31:0];
   assign R8     = s_logisimBus38[31:0];
   assign R9     = s_logisimBus22[31:0];

   /*******************************************************************************
   ** Here all in-lined components are defined                                   **
   *******************************************************************************/

   // Constant
   assign  s_logisimBus52[31:0]  =  32'h00000000;


   // Constant
   assign  s_logisimBus41[31:0]  =  32'h00000000;


   // Constant
   assign  s_logisimBus67[31:0]  =  32'h00000000;


   /*******************************************************************************
   ** Here all normal components are defined                                     **
   *******************************************************************************/
   AND_GATE #(.BubblesMask(2'b00))
      GATES_1 (.input1(s_logisimNet21),
               .input2(s_logisimNet51),
               .result(s_logisimNet74));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_2 (.input1(s_logisimNet21),
               .input2(s_logisimNet25),
               .result(s_logisimNet75));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_3 (.input1(s_logisimNet21),
               .input2(s_logisimNet20),
               .result(s_logisimNet76));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_4 (.input1(s_logisimNet21),
               .input2(s_logisimNet5),
               .result(s_logisimNet77));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_5 (.input1(s_logisimNet21),
               .input2(s_logisimNet18),
               .result(s_logisimNet78));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_6 (.input1(s_logisimNet21),
               .input2(s_logisimNet9),
               .result(s_logisimNet79));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_7 (.input1(s_logisimNet21),
               .input2(s_logisimNet15),
               .result(s_logisimNet80));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_8 (.input1(s_logisimNet21),
               .input2(s_logisimNet34),
               .result(s_logisimNet81));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_9 (.input1(s_logisimNet6),
               .input2(s_logisimNet74),
               .result(s_logisimNet113));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_10 (.input1(s_logisimNet6),
                .input2(s_logisimNet75),
                .result(s_logisimNet106));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_11 (.input1(s_logisimNet6),
                .input2(s_logisimNet76),
                .result(s_logisimNet107));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_12 (.input1(s_logisimNet6),
                .input2(s_logisimNet77),
                .result(s_logisimNet108));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_13 (.input1(s_logisimNet6),
                .input2(s_logisimNet78),
                .result(s_logisimNet109));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_14 (.input1(s_logisimNet6),
                .input2(s_logisimNet79),
                .result(s_logisimNet110));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_15 (.input1(s_logisimNet6),
                .input2(s_logisimNet80),
                .result(s_logisimNet111));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_16 (.input1(s_logisimNet6),
                .input2(s_logisimNet81),
                .result(s_logisimNet112));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_17 (.input1(s_logisimNet64),
                .input2(s_logisimNet97),
                .result(s_logisimNet114));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_18 (.input1(s_logisimNet11),
                .input2(s_logisimNet51),
                .result(s_logisimNet82));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_19 (.input1(s_logisimNet11),
                .input2(s_logisimNet25),
                .result(s_logisimNet83));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_20 (.input1(s_logisimNet11),
                .input2(s_logisimNet20),
                .result(s_logisimNet84));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_21 (.input1(s_logisimNet11),
                .input2(s_logisimNet5),
                .result(s_logisimNet85));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_22 (.input1(s_logisimNet11),
                .input2(s_logisimNet18),
                .result(s_logisimNet86));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_23 (.input1(s_logisimNet11),
                .input2(s_logisimNet9),
                .result(s_logisimNet87));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_24 (.input1(s_logisimNet11),
                .input2(s_logisimNet15),
                .result(s_logisimNet88));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_25 (.input1(s_logisimNet11),
                .input2(s_logisimNet34),
                .result(s_logisimNet89));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_26 (.input1(s_logisimNet6),
                .input2(s_logisimNet82),
                .result(s_logisimNet122));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_27 (.input1(s_logisimNet6),
                .input2(s_logisimNet83),
                .result(s_logisimNet115));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_28 (.input1(s_logisimNet6),
                .input2(s_logisimNet84),
                .result(s_logisimNet116));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_29 (.input1(s_logisimNet6),
                .input2(s_logisimNet85),
                .result(s_logisimNet117));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_30 (.input1(s_logisimNet6),
                .input2(s_logisimNet86),
                .result(s_logisimNet118));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_31 (.input1(s_logisimNet6),
                .input2(s_logisimNet87),
                .result(s_logisimNet119));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_32 (.input1(s_logisimNet6),
                .input2(s_logisimNet88),
                .result(s_logisimNet120));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_33 (.input1(s_logisimNet6),
                .input2(s_logisimNet89),
                .result(s_logisimNet121));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_34 (.input1(s_logisimNet13),
                .input2(s_logisimNet51),
                .result(s_logisimNet90));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_35 (.input1(s_logisimNet13),
                .input2(s_logisimNet25),
                .result(s_logisimNet91));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_36 (.input1(s_logisimNet13),
                .input2(s_logisimNet20),
                .result(s_logisimNet92));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_37 (.input1(s_logisimNet13),
                .input2(s_logisimNet5),
                .result(s_logisimNet93));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_38 (.input1(s_logisimNet13),
                .input2(s_logisimNet18),
                .result(s_logisimNet94));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_39 (.input1(s_logisimNet13),
                .input2(s_logisimNet15),
                .result(s_logisimNet95));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_40 (.input1(s_logisimNet13),
                .input2(s_logisimNet34),
                .result(s_logisimNet96));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_41 (.input1(s_logisimNet6),
                .input2(s_logisimNet90),
                .result(s_logisimNet129));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_42 (.input1(s_logisimNet6),
                .input2(s_logisimNet91),
                .result(s_logisimNet123));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_43 (.input1(s_logisimNet6),
                .input2(s_logisimNet92),
                .result(s_logisimNet124));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_44 (.input1(s_logisimNet6),
                .input2(s_logisimNet93),
                .result(s_logisimNet125));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_45 (.input1(s_logisimNet6),
                .input2(s_logisimNet94),
                .result(s_logisimNet126));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_46 (.input1(s_logisimNet6),
                .input2(s_logisimNet95),
                .result(s_logisimNet127));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_47 (.input1(s_logisimNet6),
                .input2(s_logisimNet96),
                .result(s_logisimNet128));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_48 (.input1(s_logisimNet30),
                .input2(s_logisimNet51),
                .result(s_logisimNet98));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_49 (.input1(s_logisimNet30),
                .input2(s_logisimNet25),
                .result(s_logisimNet99));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_50 (.input1(s_logisimNet30),
                .input2(s_logisimNet20),
                .result(s_logisimNet100));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_51 (.input1(s_logisimNet30),
                .input2(s_logisimNet5),
                .result(s_logisimNet101));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_52 (.input1(s_logisimNet30),
                .input2(s_logisimNet18),
                .result(s_logisimNet102));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_53 (.input1(s_logisimNet30),
                .input2(s_logisimNet9),
                .result(s_logisimNet103));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_54 (.input1(s_logisimNet30),
                .input2(s_logisimNet15),
                .result(s_logisimNet104));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_55 (.input1(s_logisimNet30),
                .input2(s_logisimNet34),
                .result(s_logisimNet105));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_56 (.input1(s_logisimNet16),
                .input2(s_logisimNet66),
                .result(s_logisimNet97));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_57 (.input1(s_logisimNet6),
                .input2(s_logisimNet98),
                .result(s_logisimNet137));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_58 (.input1(s_logisimNet6),
                .input2(s_logisimNet99),
                .result(s_logisimNet130));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_59 (.input1(s_logisimNet6),
                .input2(s_logisimNet100),
                .result(s_logisimNet131));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_60 (.input1(s_logisimNet6),
                .input2(s_logisimNet101),
                .result(s_logisimNet132));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_61 (.input1(s_logisimNet6),
                .input2(s_logisimNet102),
                .result(s_logisimNet133));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_62 (.input1(s_logisimNet6),
                .input2(s_logisimNet103),
                .result(s_logisimNet134));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_63 (.input1(s_logisimNet6),
                .input2(s_logisimNet104),
                .result(s_logisimNet135));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_64 (.input1(s_logisimNet6),
                .input2(s_logisimNet105),
                .result(s_logisimNet136));

   Multiplexer_bus_8 #(.nrOfBits(32))
      PLEXERS_65 (.enable(1'b1),
                  .muxIn_0(s_logisimBus43[31:0]),
                  .muxIn_1(s_logisimBus12[31:0]),
                  .muxIn_2(s_logisimBus22[31:0]),
                  .muxIn_3(s_logisimBus24[31:0]),
                  .muxIn_4(s_logisimBus32[31:0]),
                  .muxIn_5(s_logisimBus42[31:0]),
                  .muxIn_6(s_logisimBus33[31:0]),
                  .muxIn_7(s_logisimBus35[31:0]),
                  .muxOut(s_logisimBus47[31:0]),
                  .sel(s_logisimBus55[4:2]));

   Multiplexer_bus_8 #(.nrOfBits(32))
      PLEXERS_66 (.enable(1'b1),
                  .muxIn_0(s_logisimBus43[31:0]),
                  .muxIn_1(s_logisimBus12[31:0]),
                  .muxIn_2(s_logisimBus22[31:0]),
                  .muxIn_3(s_logisimBus24[31:0]),
                  .muxIn_4(s_logisimBus32[31:0]),
                  .muxIn_5(s_logisimBus42[31:0]),
                  .muxIn_6(s_logisimBus33[31:0]),
                  .muxIn_7(s_logisimBus35[31:0]),
                  .muxOut(s_logisimBus72[31:0]),
                  .sel(s_logisimBus37[4:2]));

   Multiplexer_bus_8 #(.nrOfBits(32))
      PLEXERS_67 (.enable(1'b1),
                  .muxIn_0(s_logisimBus27[31:0]),
                  .muxIn_1(s_logisimBus40[31:0]),
                  .muxIn_2(s_logisimBus44[31:0]),
                  .muxIn_3(s_logisimBus45[31:0]),
                  .muxIn_4(s_logisimBus1[31:0]),
                  .muxIn_5(s_logisimBus53[31:0]),
                  .muxIn_6(s_logisimBus49[31:0]),
                  .muxIn_7(s_logisimBus50[31:0]),
                  .muxOut(s_logisimBus71[31:0]),
                  .sel(s_logisimBus55[4:2]));

   Multiplexer_bus_8 #(.nrOfBits(32))
      PLEXERS_68 (.enable(1'b1),
                  .muxIn_0(s_logisimBus27[31:0]),
                  .muxIn_1(s_logisimBus40[31:0]),
                  .muxIn_2(s_logisimBus44[31:0]),
                  .muxIn_3(s_logisimBus45[31:0]),
                  .muxIn_4(s_logisimBus1[31:0]),
                  .muxIn_5(s_logisimBus53[31:0]),
                  .muxIn_6(s_logisimBus49[31:0]),
                  .muxIn_7(s_logisimBus50[31:0]),
                  .muxOut(s_logisimBus68[31:0]),
                  .sel(s_logisimBus37[4:2]));

   Multiplexer_bus_8 #(.nrOfBits(32))
      PLEXERS_69 (.enable(1'b1),
                  .muxIn_0(s_logisimBus46[31:0]),
                  .muxIn_1(s_logisimBus23[31:0]),
                  .muxIn_2(s_logisimBus54[31:0]),
                  .muxIn_3(s_logisimBus56[31:0]),
                  .muxIn_4(s_logisimBus31[31:0]),
                  .muxIn_5(s_logisimBus62[31:0]),
                  .muxIn_6(s_logisimBus28[31:0]),
                  .muxIn_7(s_logisimBus59[31:0]),
                  .muxOut(s_logisimBus39[31:0]),
                  .sel(s_logisimBus55[4:2]));

   Multiplexer_bus_8 #(.nrOfBits(32))
      PLEXERS_70 (.enable(1'b1),
                  .muxIn_0(s_logisimBus46[31:0]),
                  .muxIn_1(s_logisimBus23[31:0]),
                  .muxIn_2(s_logisimBus54[31:0]),
                  .muxIn_3(s_logisimBus56[31:0]),
                  .muxIn_4(s_logisimBus31[31:0]),
                  .muxIn_5(s_logisimBus62[31:0]),
                  .muxIn_6(s_logisimBus28[31:0]),
                  .muxIn_7(s_logisimBus59[31:0]),
                  .muxOut(s_logisimBus8[31:0]),
                  .sel(s_logisimBus37[4:2]));

   Multiplexer_bus_4 #(.nrOfBits(32))
      PLEXERS_71 (.enable(1'b1),
                  .muxIn_0(s_logisimBus10[31:0]),
                  .muxIn_1(s_logisimBus72[31:0]),
                  .muxIn_2(s_logisimBus68[31:0]),
                  .muxIn_3(s_logisimBus8[31:0]),
                  .muxOut(s_logisimBus70[31:0]),
                  .sel(s_logisimBus37[1:0]));

   Multiplexer_bus_4 #(.nrOfBits(32))
      PLEXERS_72 (.enable(1'b1),
                  .muxIn_0(s_logisimBus61[31:0]),
                  .muxIn_1(s_logisimBus47[31:0]),
                  .muxIn_2(s_logisimBus71[31:0]),
                  .muxIn_3(s_logisimBus39[31:0]),
                  .muxOut(s_logisimBus63[31:0]),
                  .sel(s_logisimBus55[1:0]));

   Decoder_8   PLEXERS_73 (.decoderOut_0(s_logisimNet9),
                           .decoderOut_1(s_logisimNet15),
                           .decoderOut_2(s_logisimNet34),
                           .decoderOut_3(s_logisimNet51),
                           .decoderOut_4(s_logisimNet25),
                           .decoderOut_5(s_logisimNet20),
                           .decoderOut_6(s_logisimNet5),
                           .decoderOut_7(s_logisimNet18),
                           .enable(1'b1),
                           .sel(s_logisimBus17[4:2]));

   Decoder_4   PLEXERS_74 (.decoderOut_0(s_logisimNet13),
                           .decoderOut_1(s_logisimNet30),
                           .decoderOut_2(s_logisimNet21),
                           .decoderOut_3(s_logisimNet11),
                           .enable(1'b1),
                           .sel(s_logisimBus17[1:0]));

   Multiplexer_bus_2 #(.nrOfBits(32))
      PLEXERS_75 (.enable(1'b1),
                  .muxIn_0(s_logisimBus73[31:0]),
                  .muxIn_1(s_logisimBus52[31:0]),
                  .muxOut(s_logisimBus0[31:0]),
                  .sel(s_logisimNet6));

   Multiplexer_bus_8 #(.nrOfBits(32))
      PLEXERS_76 (.enable(1'b1),
                  .muxIn_0(s_logisimBus41[31:0]),
                  .muxIn_1(s_logisimBus58[31:0]),
                  .muxIn_2(s_logisimBus38[31:0]),
                  .muxIn_3(s_logisimBus14[31:0]),
                  .muxIn_4(s_logisimBus2[31:0]),
                  .muxIn_5(s_logisimBus19[31:0]),
                  .muxIn_6(s_logisimBus7[31:0]),
                  .muxIn_7(s_logisimBus29[31:0]),
                  .muxOut(s_logisimBus61[31:0]),
                  .sel(s_logisimBus55[4:2]));

   Multiplexer_bus_8 #(.nrOfBits(32))
      PLEXERS_77 (.enable(1'b1),
                  .muxIn_0(s_logisimBus67[31:0]),
                  .muxIn_1(s_logisimBus58[31:0]),
                  .muxIn_2(s_logisimBus38[31:0]),
                  .muxIn_3(s_logisimBus14[31:0]),
                  .muxIn_4(s_logisimBus2[31:0]),
                  .muxIn_5(s_logisimBus19[31:0]),
                  .muxIn_6(s_logisimBus7[31:0]),
                  .muxIn_7(s_logisimBus29[31:0]),
                  .muxOut(s_logisimBus10[31:0]),
                  .sel(s_logisimBus37[4:2]));

   REGISTER_FLIP_FLOP #(.invertClock(0),
                        .nrOfBits(32))
      MEMORY_78 (.clock(s_logisimNet3),
                 .clockEnable(s_logisimNet106),
                 .d(s_logisimBus0[31:0]),
                 .q(s_logisimBus1[31:0]),
                 .reset(1'b0),
                 .tick(1'b1));

   REGISTER_FLIP_FLOP #(.invertClock(0),
                        .nrOfBits(32))
      MEMORY_79 (.clock(s_logisimNet3),
                 .clockEnable(s_logisimNet107),
                 .d(s_logisimBus0[31:0]),
                 .q(s_logisimBus53[31:0]),
                 .reset(1'b0),
                 .tick(1'b1));

   REGISTER_FLIP_FLOP #(.invertClock(0),
                        .nrOfBits(32))
      MEMORY_80 (.clock(s_logisimNet3),
                 .clockEnable(s_logisimNet108),
                 .d(s_logisimBus0[31:0]),
                 .q(s_logisimBus49[31:0]),
                 .reset(1'b0),
                 .tick(1'b1));

   REGISTER_FLIP_FLOP #(.invertClock(0),
                        .nrOfBits(32))
      MEMORY_81 (.clock(s_logisimNet3),
                 .clockEnable(s_logisimNet109),
                 .d(s_logisimBus0[31:0]),
                 .q(s_logisimBus50[31:0]),
                 .reset(1'b0),
                 .tick(1'b1));

   REGISTER_FLIP_FLOP #(.invertClock(0),
                        .nrOfBits(32))
      MEMORY_82 (.clock(s_logisimNet3),
                 .clockEnable(s_logisimNet110),
                 .d(s_logisimBus0[31:0]),
                 .q(s_logisimBus27[31:0]),
                 .reset(1'b0),
                 .tick(1'b1));

   REGISTER_FLIP_FLOP #(.invertClock(0),
                        .nrOfBits(32))
      MEMORY_83 (.clock(s_logisimNet3),
                 .clockEnable(s_logisimNet111),
                 .d(s_logisimBus0[31:0]),
                 .q(s_logisimBus40[31:0]),
                 .reset(1'b0),
                 .tick(1'b1));

   REGISTER_FLIP_FLOP #(.invertClock(0),
                        .nrOfBits(32))
      MEMORY_84 (.clock(s_logisimNet3),
                 .clockEnable(s_logisimNet112),
                 .d(s_logisimBus0[31:0]),
                 .q(s_logisimBus44[31:0]),
                 .reset(1'b0),
                 .tick(1'b1));

   REGISTER_FLIP_FLOP #(.invertClock(0),
                        .nrOfBits(32))
      MEMORY_85 (.clock(s_logisimNet3),
                 .clockEnable(s_logisimNet113),
                 .d(s_logisimBus0[31:0]),
                 .q(s_logisimBus45[31:0]),
                 .reset(1'b0),
                 .tick(1'b1));

   REGISTER_FLIP_FLOP #(.invertClock(0),
                        .nrOfBits(32))
      MEMORY_86 (.clock(s_logisimNet26),
                 .clockEnable(s_logisimNet114),
                 .d(s_logisimBus36[31:0]),
                 .q(),
                 .reset(1'b0),
                 .tick(1'b1));

   REGISTER_FLIP_FLOP #(.invertClock(0),
                        .nrOfBits(32))
      MEMORY_87 (.clock(s_logisimNet3),
                 .clockEnable(s_logisimNet115),
                 .d(s_logisimBus0[31:0]),
                 .q(s_logisimBus31[31:0]),
                 .reset(1'b0),
                 .tick(1'b1));

   REGISTER_FLIP_FLOP #(.invertClock(0),
                        .nrOfBits(32))
      MEMORY_88 (.clock(s_logisimNet3),
                 .clockEnable(s_logisimNet116),
                 .d(s_logisimBus0[31:0]),
                 .q(s_logisimBus62[31:0]),
                 .reset(1'b0),
                 .tick(1'b1));

   REGISTER_FLIP_FLOP #(.invertClock(0),
                        .nrOfBits(32))
      MEMORY_89 (.clock(s_logisimNet3),
                 .clockEnable(s_logisimNet117),
                 .d(s_logisimBus0[31:0]),
                 .q(s_logisimBus28[31:0]),
                 .reset(1'b0),
                 .tick(1'b1));

   REGISTER_FLIP_FLOP #(.invertClock(0),
                        .nrOfBits(32))
      MEMORY_90 (.clock(s_logisimNet3),
                 .clockEnable(s_logisimNet118),
                 .d(s_logisimBus0[31:0]),
                 .q(s_logisimBus59[31:0]),
                 .reset(1'b0),
                 .tick(1'b1));

   REGISTER_FLIP_FLOP #(.invertClock(0),
                        .nrOfBits(32))
      MEMORY_91 (.clock(s_logisimNet3),
                 .clockEnable(s_logisimNet119),
                 .d(s_logisimBus0[31:0]),
                 .q(s_logisimBus46[31:0]),
                 .reset(1'b0),
                 .tick(1'b1));

   REGISTER_FLIP_FLOP #(.invertClock(0),
                        .nrOfBits(32))
      MEMORY_92 (.clock(s_logisimNet3),
                 .clockEnable(s_logisimNet120),
                 .d(s_logisimBus0[31:0]),
                 .q(s_logisimBus23[31:0]),
                 .reset(1'b0),
                 .tick(1'b1));

   REGISTER_FLIP_FLOP #(.invertClock(0),
                        .nrOfBits(32))
      MEMORY_93 (.clock(s_logisimNet3),
                 .clockEnable(s_logisimNet121),
                 .d(s_logisimBus0[31:0]),
                 .q(s_logisimBus54[31:0]),
                 .reset(1'b0),
                 .tick(1'b1));

   REGISTER_FLIP_FLOP #(.invertClock(0),
                        .nrOfBits(32))
      MEMORY_94 (.clock(s_logisimNet3),
                 .clockEnable(s_logisimNet122),
                 .d(s_logisimBus0[31:0]),
                 .q(s_logisimBus56[31:0]),
                 .reset(1'b0),
                 .tick(1'b1));

   REGISTER_FLIP_FLOP #(.invertClock(0),
                        .nrOfBits(32))
      MEMORY_95 (.clock(s_logisimNet3),
                 .clockEnable(s_logisimNet123),
                 .d(s_logisimBus0[31:0]),
                 .q(s_logisimBus2[31:0]),
                 .reset(1'b0),
                 .tick(1'b1));

   REGISTER_FLIP_FLOP #(.invertClock(0),
                        .nrOfBits(32))
      MEMORY_96 (.clock(s_logisimNet3),
                 .clockEnable(s_logisimNet124),
                 .d(s_logisimBus0[31:0]),
                 .q(s_logisimBus19[31:0]),
                 .reset(1'b0),
                 .tick(1'b1));

   REGISTER_FLIP_FLOP #(.invertClock(0),
                        .nrOfBits(32))
      MEMORY_97 (.clock(s_logisimNet3),
                 .clockEnable(s_logisimNet125),
                 .d(s_logisimBus0[31:0]),
                 .q(s_logisimBus7[31:0]),
                 .reset(1'b0),
                 .tick(1'b1));

   REGISTER_FLIP_FLOP #(.invertClock(0),
                        .nrOfBits(32))
      MEMORY_98 (.clock(s_logisimNet3),
                 .clockEnable(s_logisimNet126),
                 .d(s_logisimBus0[31:0]),
                 .q(s_logisimBus29[31:0]),
                 .reset(1'b0),
                 .tick(1'b1));

   REGISTER_FLIP_FLOP #(.invertClock(0),
                        .nrOfBits(32))
      MEMORY_99 (.clock(s_logisimNet3),
                 .clockEnable(s_logisimNet127),
                 .d(s_logisimBus0[31:0]),
                 .q(s_logisimBus58[31:0]),
                 .reset(1'b0),
                 .tick(1'b1));

   REGISTER_FLIP_FLOP #(.invertClock(0),
                        .nrOfBits(32))
      MEMORY_100 (.clock(s_logisimNet3),
                  .clockEnable(s_logisimNet128),
                  .d(s_logisimBus0[31:0]),
                  .q(s_logisimBus38[31:0]),
                  .reset(1'b0),
                  .tick(1'b1));

   REGISTER_FLIP_FLOP #(.invertClock(0),
                        .nrOfBits(32))
      MEMORY_101 (.clock(s_logisimNet3),
                  .clockEnable(s_logisimNet129),
                  .d(s_logisimBus0[31:0]),
                  .q(s_logisimBus14[31:0]),
                  .reset(1'b0),
                  .tick(1'b1));

   REGISTER_FLIP_FLOP #(.invertClock(0),
                        .nrOfBits(32))
      MEMORY_102 (.clock(s_logisimNet3),
                  .clockEnable(s_logisimNet130),
                  .d(s_logisimBus0[31:0]),
                  .q(s_logisimBus32[31:0]),
                  .reset(1'b0),
                  .tick(1'b1));

   REGISTER_FLIP_FLOP #(.invertClock(0),
                        .nrOfBits(32))
      MEMORY_103 (.clock(s_logisimNet3),
                  .clockEnable(s_logisimNet131),
                  .d(s_logisimBus0[31:0]),
                  .q(s_logisimBus42[31:0]),
                  .reset(1'b0),
                  .tick(1'b1));

   REGISTER_FLIP_FLOP #(.invertClock(0),
                        .nrOfBits(32))
      MEMORY_104 (.clock(s_logisimNet3),
                  .clockEnable(s_logisimNet132),
                  .d(s_logisimBus0[31:0]),
                  .q(s_logisimBus33[31:0]),
                  .reset(1'b0),
                  .tick(1'b1));

   REGISTER_FLIP_FLOP #(.invertClock(0),
                        .nrOfBits(32))
      MEMORY_105 (.clock(s_logisimNet3),
                  .clockEnable(s_logisimNet133),
                  .d(s_logisimBus0[31:0]),
                  .q(s_logisimBus35[31:0]),
                  .reset(1'b0),
                  .tick(1'b1));

   REGISTER_FLIP_FLOP #(.invertClock(0),
                        .nrOfBits(32))
      MEMORY_106 (.clock(s_logisimNet3),
                  .clockEnable(s_logisimNet134),
                  .d(s_logisimBus0[31:0]),
                  .q(s_logisimBus43[31:0]),
                  .reset(1'b0),
                  .tick(1'b1));

   REGISTER_FLIP_FLOP #(.invertClock(0),
                        .nrOfBits(32))
      MEMORY_107 (.clock(s_logisimNet3),
                  .clockEnable(s_logisimNet135),
                  .d(s_logisimBus0[31:0]),
                  .q(s_logisimBus12[31:0]),
                  .reset(1'b0),
                  .tick(1'b1));

   REGISTER_FLIP_FLOP #(.invertClock(0),
                        .nrOfBits(32))
      MEMORY_108 (.clock(s_logisimNet3),
                  .clockEnable(s_logisimNet136),
                  .d(s_logisimBus0[31:0]),
                  .q(s_logisimBus22[31:0]),
                  .reset(1'b0),
                  .tick(1'b1));

   REGISTER_FLIP_FLOP #(.invertClock(0),
                        .nrOfBits(32))
      MEMORY_109 (.clock(s_logisimNet3),
                  .clockEnable(s_logisimNet137),
                  .d(s_logisimBus0[31:0]),
                  .q(s_logisimBus24[31:0]),
                  .reset(1'b0),
                  .tick(1'b1));


endmodule
