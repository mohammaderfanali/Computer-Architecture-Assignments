/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
Control_Unit
**
**
**
*****************************************************************************/
module
Control_Unit(
Opcode,
aluop,
beq,
bne,
funct,
is_div,
is_jal,
is_jr,
is_mul,
jump,
lo_or_hi,
mem_to_reg,
mem_write,
mf,
reg_write,
regdst,
sll_control,
slti,
source_2
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[5:0]
Opcode;
input
[5:0]
funct;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
[3:0]
aluop;
output
beq;
output
bne;
output
is_div;
output
is_jal;
output
is_jr;
output
is_mul;
output
jump;
output
lo_or_hi;
output
mem_to_reg;
output
mem_write;
output
mf;
output
reg_write;
output
regdst;
output
sll_control;
output
slti;
output
source_2;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[5:0]
s_logisimBus1;
wire
[5:0]
s_logisimBus11;
wire
[5:0]
s_logisimBus12;
wire
[5:0]
s_logisimBus13;
wire
[5:0]
s_logisimBus14;
wire
[5:0]
s_logisimBus24;
wire
[5:0]
s_logisimBus31;
wire
[5:0]
s_logisimBus36;
wire
[5:0]
s_logisimBus37;
wire
[3:0]
s_logisimBus38;
wire
[5:0]
s_logisimBus42;
wire
[5:0]
s_logisimBus46;
wire
[5:0]
s_logisimBus48;
wire
[5:0]
s_logisimBus49;
wire
[5:0]
s_logisimBus50;
wire
[5:0]
s_logisimBus51;
wire
[5:0]
s_logisimBus52;
wire
[5:0]
s_logisimBus53;
wire
s_logisimNet0;
wire
s_logisimNet10;
wire
s_logisimNet15;
wire
s_logisimNet16;
wire
s_logisimNet17;
wire
s_logisimNet18;
wire
s_logisimNet19;
wire
s_logisimNet2;
wire
s_logisimNet20;
wire
s_logisimNet21;
wire
s_logisimNet22;
wire
s_logisimNet23;
wire
s_logisimNet25;
wire
s_logisimNet26;
wire
s_logisimNet27;
wire
s_logisimNet28;
wire
s_logisimNet29;
wire
s_logisimNet3;
wire
s_logisimNet30;
wire
s_logisimNet32;
wire
s_logisimNet33;
wire
s_logisimNet34;
wire
s_logisimNet35;
wire
s_logisimNet39;
wire
s_logisimNet4;
wire
s_logisimNet40;
wire
s_logisimNet41;
wire
s_logisimNet43;
wire
s_logisimNet44;
wire
s_logisimNet45;
wire
s_logisimNet47;
wire
s_logisimNet5;
wire
s_logisimNet54;
wire
s_logisimNet55;
wire
s_logisimNet56;
wire
s_logisimNet57;
wire
s_logisimNet58;
wire
s_logisimNet59;
wire
s_logisimNet6;
wire
s_logisimNet60;
wire
s_logisimNet61;
wire
s_logisimNet7;
wire
s_logisimNet8;
wire
s_logisimNet9;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus13[5:0]
=
funct;
assign
s_logisimBus1[5:0]
=
Opcode;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
aluop
=
s_logisimBus38[3:0];
assign
beq
=
s_logisimNet40;
assign
bne
=
s_logisimNet23;
assign
is_div
=
s_logisimNet6;
assign
is_jal
=
s_logisimNet56;
assign
is_jr
=
s_logisimNet3;
assign
is_mul
=
s_logisimNet58;
assign
jump
=
s_logisimNet60;
assign
lo_or_hi
=
s_logisimBus13[1];
assign
mem_to_reg
=
s_logisimNet59;
assign
mem_write
=
s_logisimNet43;
assign
mf
=
s_logisimNet4;
assign
reg_write
=
s_logisimNet25;
assign
regdst
=
s_logisimNet26;
assign
sll_control
=
s_logisimNet29;
assign
slti
=
s_logisimNet16;
assign
source_2
=
s_logisimNet45;
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus52[5:0]
=
{2'b01,
4'hC};
assign
s_logisimBus48[5:0]
=
{2'b00,
4'h0};
assign
s_logisimBus11[5:0]
=
{2'b00,
4'h8};
assign
s_logisimBus46[5:0]
=
{2'b00,
4'h8};
assign
s_logisimBus49[5:0]
=
{2'b00,
4'h3};
assign
s_logisimBus42[5:0]
=
{2'b10,
4'h3};
assign
s_logisimBus50[5:0]
=
{2'b00,
4'hA};
assign
s_logisimBus53[5:0]
=
{2'b00,
4'h0};
assign
s_logisimBus24[5:0]
=
{2'b01,
4'hC};
assign
s_logisimBus31[5:0]
=
{2'b00,
4'h2};
assign
s_logisimBus37[5:0]
=
{2'b00,
4'h4};
assign
s_logisimBus36[5:0]
=
{2'b10,
4'hB};
assign
s_logisimBus14[5:0]
=
{2'b01,
4'hA};
assign
s_logisimBus51[5:0]
=
{2'b00,
4'h8};
assign
s_logisimBus12[5:0]
=
{2'b00,
4'h5};
assign
s_logisimNet15
=
~s_logisimBus1[3];
assign
s_logisimNet47
=
~s_logisimBus1[1];
assign
s_logisimNet32
=
~s_logisimBus1[0];
assign
s_logisimNet21
=
~s_logisimBus13[3];
assign
s_logisimNet26
=
~s_logisimNet61;
assign
s_logisimNet35
=
~s_logisimNet6;
assign
s_logisimNet22
=
~s_logisimNet8;
assign
s_logisimNet33
=
~s_logisimNet28;
assign
s_logisimNet34
=
~s_logisimNet44;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
AND_GATE_3_INPUTS
#(.BubblesMask(3'b000))
GATES_1
(.input1(s_logisimNet26),
.input2(s_logisimNet22),
.input3(s_logisimNet33),
.result(s_logisimNet45));
OR_GATE
#(.BubblesMask(2'b00))
GATES_2
(.input1(s_logisimNet5),
.input2(s_logisimNet9),
.result(s_logisimNet61));
AND_GATE_3_INPUTS
#(.BubblesMask(3'b000))
GATES_3
(.input1(s_logisimNet32),
.input2(s_logisimBus1[1]),
.input3(s_logisimNet15),
.result(s_logisimNet55));
AND_GATE_3_INPUTS
#(.BubblesMask(3'b000))
GATES_4
(.input1(s_logisimBus1[0]),
.input2(s_logisimNet47),
.input3(s_logisimBus1[2]),
.result(s_logisimNet23));
OR_GATE
#(.BubblesMask(2'b00))
GATES_5
(.input1(s_logisimNet55),
.input2(s_logisimNet56),
.result(s_logisimNet60));
AND_GATE_3_INPUTS
#(.BubblesMask(3'b000))
GATES_6
(.input1(s_logisimNet61),
.input2(s_logisimNet21),
.input3(s_logisimBus13[4]),
.result(s_logisimNet4));
OR_GATE_4_INPUTS
#(.BubblesMask(4'h0))
GATES_7
(.input1(s_logisimNet10),
.input2(s_logisimNet61),
.input3(s_logisimNet2),
.input4(s_logisimNet16),
.result(s_logisimNet20));
AND_GATE
#(.BubblesMask(2'b00))
GATES_8
(.input1(s_logisimNet61),
.input2(s_logisimNet41),
.result(s_logisimNet29));
AND_GATE
#(.BubblesMask(2'b00))
GATES_9
(.input1(s_logisimNet61),
.input2(s_logisimNet39),
.result(s_logisimNet6));
AND_GATE
#(.BubblesMask(2'b00))
GATES_10
(.input1(s_logisimNet8),
.input2(s_logisimNet18),
.result(s_logisimNet58));
AND_GATE
#(.BubblesMask(2'b00))
GATES_11
(.input1(s_logisimNet61),
.input2(s_logisimNet54),
.result(s_logisimNet3));
AND_GATE
#(.BubblesMask(2'b00))
GATES_12
(.input1(s_logisimNet20),
.input2(s_logisimNet35),
.result(s_logisimNet25));
AND_GATE
#(.BubblesMask(2'b00))
GATES_13
(.input1(s_logisimNet26),
.input2(s_logisimNet34),
.result(s_logisimNet59));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_14
(.aEqualsB(s_logisimNet5),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus52[5:0]),
.dataB(s_logisimBus1[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_15
(.aEqualsB(s_logisimNet9),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus48[5:0]),
.dataB(s_logisimBus1[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(1))
ARITH_16
(.aEqualsB(s_logisimNet54),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus13[5:0]),
.dataB(s_logisimBus11[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_17
(.aEqualsB(s_logisimNet10),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus46[5:0]),
.dataB(s_logisimBus1[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_18
(.aEqualsB(s_logisimNet56),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus49[5:0]),
.dataB(s_logisimBus1[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_19
(.aEqualsB(s_logisimNet2),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus1[5:0]),
.dataB(s_logisimBus42[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_20
(.aEqualsB(s_logisimNet16),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus1[5:0]),
.dataB(s_logisimBus50[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_21
(.aEqualsB(s_logisimNet41),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus53[5:0]),
.dataB(s_logisimBus13[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_22
(.aEqualsB(),
.aGreaterThanB(),
.aLessThanB(),
.dataA(6'd0),
.dataB(6'd0));
Comparator
#(.nrOfBits(6),
.twosComplement(1))
ARITH_23
(.aEqualsB(s_logisimNet8),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus1[5:0]),
.dataB(s_logisimBus24[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(1))
ARITH_24
(.aEqualsB(s_logisimNet18),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus13[5:0]),
.dataB(s_logisimBus31[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(1))
ARITH_25
(.aEqualsB(s_logisimNet40),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus1[5:0]),
.dataB(s_logisimBus37[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_26
(.aEqualsB(s_logisimNet39),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus13[5:0]),
.dataB(s_logisimBus14[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_27
(.aEqualsB(s_logisimNet43),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus36[5:0]),
.dataB(s_logisimBus1[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_28
(.aEqualsB(s_logisimNet28),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus12[5:0]),
.dataB(s_logisimBus1[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_29
(.aEqualsB(s_logisimNet44),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus51[5:0]),
.dataB(s_logisimBus1[5:0]));
/*******************************************************************************
**
Here
all
sub-circuits
are
defined
**
*******************************************************************************/
Control_Alu
alu_controler
(.Opcode(s_logisimBus1[5:0]),
.aluop(s_logisimBus38[3:0]),
.funct(s_logisimBus13[5:0]));
endmodule