/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
main
**
**
**
*****************************************************************************/
module
main(
InstDone,
Jen,
Jin,
Jout,
R1,
R10,
R11,
R12,
R13,
R14,
R15,
R16,
R17,
R18,
R19,
R2,
R20,
R21,
R22,
R23,
R24,
R25,
R26,
R27,
R28,
R29,
R3,
R30,
R31,
R4,
R5,
R6,
R7,
R8,
R9,
clk,
rst
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
Jen;
input
[31:0]
Jin;
input
clk;
input
rst;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
InstDone;
output
[31:0]
Jout;
output
[31:0]
R1;
output
[31:0]
R10;
output
[31:0]
R11;
output
[31:0]
R12;
output
[31:0]
R13;
output
[31:0]
R14;
output
[31:0]
R15;
output
[31:0]
R16;
output
[31:0]
R17;
output
[31:0]
R18;
output
[31:0]
R19;
output
[31:0]
R2;
output
[31:0]
R20;
output
[31:0]
R21;
output
[31:0]
R22;
output
[31:0]
R23;
output
[31:0]
R24;
output
[31:0]
R25;
output
[31:0]
R26;
output
[31:0]
R27;
output
[31:0]
R28;
output
[31:0]
R29;
output
[31:0]
R3;
output
[31:0]
R30;
output
[31:0]
R31;
output
[31:0]
R4;
output
[31:0]
R5;
output
[31:0]
R6;
output
[31:0]
R7;
output
[31:0]
R8;
output
[31:0]
R9;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[31:0]
s_logisimBus0;
wire
[31:0]
s_logisimBus1;
wire
[8:0]
s_logisimBus10;
wire
[31:0]
s_logisimBus100;
wire
[31:0]
s_logisimBus101;
wire
[31:0]
s_logisimBus102;
wire
[31:0]
s_logisimBus103;
wire
[31:0]
s_logisimBus104;
wire
[31:0]
s_logisimBus105;
wire
[31:0]
s_logisimBus106;
wire
[31:0]
s_logisimBus107;
wire
[31:0]
s_logisimBus108;
wire
[31:0]
s_logisimBus109;
wire
[31:0]
s_logisimBus11;
wire
[31:0]
s_logisimBus110;
wire
[31:0]
s_logisimBus111;
wire
[31:0]
s_logisimBus112;
wire
[31:0]
s_logisimBus113;
wire
[31:0]
s_logisimBus114;
wire
[31:0]
s_logisimBus115;
wire
[31:0]
s_logisimBus116;
wire
[31:0]
s_logisimBus117;
wire
[31:0]
s_logisimBus118;
wire
[31:0]
s_logisimBus119;
wire
[31:0]
s_logisimBus12;
wire
[31:0]
s_logisimBus120;
wire
[31:0]
s_logisimBus121;
wire
[31:0]
s_logisimBus122;
wire
[31:0]
s_logisimBus123;
wire
[31:0]
s_logisimBus124;
wire
[31:0]
s_logisimBus125;
wire
[31:0]
s_logisimBus126;
wire
[31:0]
s_logisimBus127;
wire
[31:0]
s_logisimBus128;
wire
[31:0]
s_logisimBus129;
wire
[8:0]
s_logisimBus13;
wire
[31:0]
s_logisimBus16;
wire
[8:0]
s_logisimBus17;
wire
[8:0]
s_logisimBus24;
wire
[31:0]
s_logisimBus26;
wire
[31:0]
s_logisimBus28;
wire
[8:0]
s_logisimBus29;
wire
[31:0]
s_logisimBus3;
wire
[8:0]
s_logisimBus30;
wire
[8:0]
s_logisimBus31;
wire
[31:0]
s_logisimBus32;
wire
[31:0]
s_logisimBus34;
wire
[4:0]
s_logisimBus37;
wire
[31:0]
s_logisimBus38;
wire
[31:0]
s_logisimBus39;
wire
[31:0]
s_logisimBus4;
wire
[31:0]
s_logisimBus41;
wire
[63:0]
s_logisimBus42;
wire
[8:0]
s_logisimBus47;
wire
[31:0]
s_logisimBus50;
wire
[31:0]
s_logisimBus52;
wire
[8:0]
s_logisimBus53;
wire
[31:0]
s_logisimBus55;
wire
[31:0]
s_logisimBus56;
wire
[63:0]
s_logisimBus57;
wire
[31:0]
s_logisimBus59;
wire
[4:0]
s_logisimBus6;
wire
[31:0]
s_logisimBus61;
wire
[4:0]
s_logisimBus64;
wire
[31:0]
s_logisimBus65;
wire
[31:0]
s_logisimBus66;
wire
[8:0]
s_logisimBus67;
wire
[31:0]
s_logisimBus69;
wire
[31:0]
s_logisimBus70;
wire
[31:0]
s_logisimBus74;
wire
[4:0]
s_logisimBus75;
wire
[31:0]
s_logisimBus76;
wire
[4:0]
s_logisimBus78;
wire
[8:0]
s_logisimBus79;
wire
[31:0]
s_logisimBus8;
wire
[31:0]
s_logisimBus83;
wire
[31:0]
s_logisimBus88;
wire
[31:0]
s_logisimBus9;
wire
[3:0]
s_logisimBus90;
wire
[31:0]
s_logisimBus99;
wire
s_logisimNet14;
wire
s_logisimNet15;
wire
s_logisimNet18;
wire
s_logisimNet19;
wire
s_logisimNet2;
wire
s_logisimNet20;
wire
s_logisimNet21;
wire
s_logisimNet22;
wire
s_logisimNet23;
wire
s_logisimNet27;
wire
s_logisimNet33;
wire
s_logisimNet35;
wire
s_logisimNet40;
wire
s_logisimNet44;
wire
s_logisimNet46;
wire
s_logisimNet48;
wire
s_logisimNet49;
wire
s_logisimNet51;
wire
s_logisimNet54;
wire
s_logisimNet58;
wire
s_logisimNet62;
wire
s_logisimNet63;
wire
s_logisimNet68;
wire
s_logisimNet71;
wire
s_logisimNet73;
wire
s_logisimNet80;
wire
s_logisimNet81;
wire
s_logisimNet82;
wire
s_logisimNet84;
wire
s_logisimNet86;
wire
s_logisimNet87;
wire
s_logisimNet89;
wire
s_logisimNet91;
wire
s_logisimNet92;
wire
s_logisimNet93;
wire
s_logisimNet94;
wire
s_logisimNet95;
wire
s_logisimNet96;
wire
s_logisimNet97;
wire
s_logisimNet98;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus41[31:0]
=
Jin;
assign
s_logisimNet35
=
Jen;
assign
s_logisimNet80
=
rst;
assign
s_logisimNet95
=
clk;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
InstDone
=
s_logisimNet54;
assign
Jout
=
s_logisimBus83[31:0];
assign
R1
=
s_logisimBus99[31:0];
assign
R10
=
s_logisimBus108[31:0];
assign
R11
=
s_logisimBus109[31:0];
assign
R12
=
s_logisimBus110[31:0];
assign
R13
=
s_logisimBus111[31:0];
assign
R14
=
s_logisimBus112[31:0];
assign
R15
=
s_logisimBus113[31:0];
assign
R16
=
s_logisimBus114[31:0];
assign
R17
=
s_logisimBus115[31:0];
assign
R18
=
s_logisimBus116[31:0];
assign
R19
=
s_logisimBus117[31:0];
assign
R2
=
s_logisimBus100[31:0];
assign
R20
=
s_logisimBus118[31:0];
assign
R21
=
s_logisimBus119[31:0];
assign
R22
=
s_logisimBus120[31:0];
assign
R23
=
s_logisimBus121[31:0];
assign
R24
=
s_logisimBus122[31:0];
assign
R25
=
s_logisimBus123[31:0];
assign
R26
=
s_logisimBus124[31:0];
assign
R27
=
s_logisimBus125[31:0];
assign
R28
=
s_logisimBus126[31:0];
assign
R29
=
s_logisimBus127[31:0];
assign
R3
=
s_logisimBus101[31:0];
assign
R30
=
s_logisimBus128[31:0];
assign
R31
=
s_logisimBus129[31:0];
assign
R4
=
s_logisimBus102[31:0];
assign
R5
=
s_logisimBus103[31:0];
assign
R6
=
s_logisimBus104[31:0];
assign
R7
=
s_logisimBus105[31:0];
assign
R8
=
s_logisimBus106[31:0];
assign
R9
=
s_logisimBus107[31:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus75[4:0]
=
{1'b1,
4'hF};
assign
s_logisimBus1[0]
=
s_logisimBus88[31];
assign
s_logisimBus1[1]
=
1'b0;
assign
s_logisimBus1[2]
=
1'b0;
assign
s_logisimBus1[3]
=
1'b0;
assign
s_logisimBus1[4]
=
1'b0;
assign
s_logisimBus1[5]
=
1'b0;
assign
s_logisimBus1[6]
=
1'b0;
assign
s_logisimBus1[7]
=
1'b0;
assign
s_logisimBus1[8]
=
1'b0;
assign
s_logisimBus1[9]
=
1'b0;
assign
s_logisimBus1[10]
=
1'b0;
assign
s_logisimBus1[11]
=
1'b0;
assign
s_logisimBus1[12]
=
1'b0;
assign
s_logisimBus1[13]
=
1'b0;
assign
s_logisimBus1[14]
=
1'b0;
assign
s_logisimBus1[15]
=
1'b0;
assign
s_logisimBus1[16]
=
1'b0;
assign
s_logisimBus1[17]
=
1'b0;
assign
s_logisimBus1[18]
=
1'b0;
assign
s_logisimBus1[19]
=
1'b0;
assign
s_logisimBus1[20]
=
1'b0;
assign
s_logisimBus1[21]
=
1'b0;
assign
s_logisimBus1[22]
=
1'b0;
assign
s_logisimBus1[23]
=
1'b0;
assign
s_logisimBus1[24]
=
1'b0;
assign
s_logisimBus1[25]
=
1'b0;
assign
s_logisimBus1[26]
=
1'b0;
assign
s_logisimBus1[27]
=
1'b0;
assign
s_logisimBus1[28]
=
1'b0;
assign
s_logisimBus1[29]
=
1'b0;
assign
s_logisimBus1[30]
=
1'b0;
assign
s_logisimBus1[31]
=
1'b0;
assign
s_logisimBus64[4:0]
=
{1'b0,
4'h0};
assign
s_logisimBus79[8:0]
=
{1'b0,
8'h01};
assign
s_logisimBus32[31:0]
=
32'h00000000;
assign
s_logisimBus34[0]
=
s_logisimBus9[0];
assign
s_logisimBus34[1]
=
s_logisimBus9[1];
assign
s_logisimBus34[2]
=
s_logisimBus9[2];
assign
s_logisimBus34[3]
=
s_logisimBus9[3];
assign
s_logisimBus34[4]
=
s_logisimBus9[4];
assign
s_logisimBus34[5]
=
s_logisimBus9[5];
assign
s_logisimBus34[6]
=
s_logisimBus9[6];
assign
s_logisimBus34[7]
=
s_logisimBus9[7];
assign
s_logisimBus34[8]
=
s_logisimBus9[8];
assign
s_logisimBus34[9]
=
s_logisimBus9[9];
assign
s_logisimBus34[10]
=
s_logisimBus9[10];
assign
s_logisimBus34[11]
=
s_logisimBus9[11];
assign
s_logisimBus34[12]
=
s_logisimBus9[12];
assign
s_logisimBus34[13]
=
s_logisimBus9[13];
assign
s_logisimBus34[14]
=
s_logisimBus9[14];
assign
s_logisimBus34[15]
=
s_logisimBus9[15];
assign
s_logisimBus34[16]
=
s_logisimBus9[15];
assign
s_logisimBus34[17]
=
s_logisimBus9[15];
assign
s_logisimBus34[18]
=
s_logisimBus9[15];
assign
s_logisimBus34[19]
=
s_logisimBus9[15];
assign
s_logisimBus34[20]
=
s_logisimBus9[15];
assign
s_logisimBus34[21]
=
s_logisimBus9[15];
assign
s_logisimBus34[22]
=
s_logisimBus9[15];
assign
s_logisimBus34[23]
=
s_logisimBus9[15];
assign
s_logisimBus34[24]
=
s_logisimBus9[15];
assign
s_logisimBus34[25]
=
s_logisimBus9[15];
assign
s_logisimBus34[26]
=
s_logisimBus9[15];
assign
s_logisimBus34[27]
=
s_logisimBus9[15];
assign
s_logisimBus34[28]
=
s_logisimBus9[15];
assign
s_logisimBus34[29]
=
s_logisimBus9[15];
assign
s_logisimBus34[30]
=
s_logisimBus9[15];
assign
s_logisimBus34[31]
=
s_logisimBus9[15];
assign
s_logisimBus8[0]
=
s_logisimBus9[6];
assign
s_logisimBus8[1]
=
s_logisimBus9[7];
assign
s_logisimBus8[2]
=
s_logisimBus9[8];
assign
s_logisimBus8[3]
=
s_logisimBus9[9];
assign
s_logisimBus8[4]
=
s_logisimBus9[10];
assign
s_logisimBus8[5]
=
s_logisimBus9[10];
assign
s_logisimBus8[6]
=
s_logisimBus9[10];
assign
s_logisimBus8[7]
=
s_logisimBus9[10];
assign
s_logisimBus8[8]
=
s_logisimBus9[10];
assign
s_logisimBus8[9]
=
s_logisimBus9[10];
assign
s_logisimBus8[10]
=
s_logisimBus9[10];
assign
s_logisimBus8[11]
=
s_logisimBus9[10];
assign
s_logisimBus8[12]
=
s_logisimBus9[10];
assign
s_logisimBus8[13]
=
s_logisimBus9[10];
assign
s_logisimBus8[14]
=
s_logisimBus9[10];
assign
s_logisimBus8[15]
=
s_logisimBus9[10];
assign
s_logisimBus8[16]
=
s_logisimBus9[10];
assign
s_logisimBus8[17]
=
s_logisimBus9[10];
assign
s_logisimBus8[18]
=
s_logisimBus9[10];
assign
s_logisimBus8[19]
=
s_logisimBus9[10];
assign
s_logisimBus8[20]
=
s_logisimBus9[10];
assign
s_logisimBus8[21]
=
s_logisimBus9[10];
assign
s_logisimBus8[22]
=
s_logisimBus9[10];
assign
s_logisimBus8[23]
=
s_logisimBus9[10];
assign
s_logisimBus8[24]
=
s_logisimBus9[10];
assign
s_logisimBus8[25]
=
s_logisimBus9[10];
assign
s_logisimBus8[26]
=
s_logisimBus9[10];
assign
s_logisimBus8[27]
=
s_logisimBus9[10];
assign
s_logisimBus8[28]
=
s_logisimBus9[10];
assign
s_logisimBus8[29]
=
s_logisimBus9[10];
assign
s_logisimBus8[30]
=
s_logisimBus9[10];
assign
s_logisimBus8[31]
=
s_logisimBus9[10];
assign
s_logisimNet19
=
1'b0;
assign
s_logisimBus4[0]
=
s_logisimBus17[0];
assign
s_logisimBus4[1]
=
s_logisimBus17[1];
assign
s_logisimBus4[2]
=
s_logisimBus17[2];
assign
s_logisimBus4[3]
=
s_logisimBus17[3];
assign
s_logisimBus4[4]
=
s_logisimBus17[4];
assign
s_logisimBus4[5]
=
s_logisimBus17[5];
assign
s_logisimBus4[6]
=
s_logisimBus17[6];
assign
s_logisimBus4[7]
=
s_logisimBus17[7];
assign
s_logisimBus4[8]
=
s_logisimBus17[8];
assign
s_logisimBus4[9]
=
1'b0;
assign
s_logisimBus4[10]
=
1'b0;
assign
s_logisimBus4[11]
=
1'b0;
assign
s_logisimBus4[12]
=
1'b0;
assign
s_logisimBus4[13]
=
1'b0;
assign
s_logisimBus4[14]
=
1'b0;
assign
s_logisimBus4[15]
=
1'b0;
assign
s_logisimBus4[16]
=
1'b0;
assign
s_logisimBus4[17]
=
1'b0;
assign
s_logisimBus4[18]
=
1'b0;
assign
s_logisimBus4[19]
=
1'b0;
assign
s_logisimBus4[20]
=
1'b0;
assign
s_logisimBus4[21]
=
1'b0;
assign
s_logisimBus4[22]
=
1'b0;
assign
s_logisimBus4[23]
=
1'b0;
assign
s_logisimBus4[24]
=
1'b0;
assign
s_logisimBus4[25]
=
1'b0;
assign
s_logisimBus4[26]
=
1'b0;
assign
s_logisimBus4[27]
=
1'b0;
assign
s_logisimBus4[28]
=
1'b0;
assign
s_logisimBus4[29]
=
1'b0;
assign
s_logisimBus4[30]
=
1'b0;
assign
s_logisimBus4[31]
=
1'b0;
assign
s_logisimBus42[0]
=
s_logisimBus88[0];
assign
s_logisimBus42[1]
=
s_logisimBus88[1];
assign
s_logisimBus42[2]
=
s_logisimBus88[2];
assign
s_logisimBus42[3]
=
s_logisimBus88[3];
assign
s_logisimBus42[4]
=
s_logisimBus88[4];
assign
s_logisimBus42[5]
=
s_logisimBus88[5];
assign
s_logisimBus42[6]
=
s_logisimBus88[6];
assign
s_logisimBus42[7]
=
s_logisimBus88[7];
assign
s_logisimBus42[8]
=
s_logisimBus88[8];
assign
s_logisimBus42[9]
=
s_logisimBus88[9];
assign
s_logisimBus42[10]
=
s_logisimBus88[10];
assign
s_logisimBus42[11]
=
s_logisimBus88[11];
assign
s_logisimBus42[12]
=
s_logisimBus88[12];
assign
s_logisimBus42[13]
=
s_logisimBus88[13];
assign
s_logisimBus42[14]
=
s_logisimBus88[14];
assign
s_logisimBus42[15]
=
s_logisimBus88[15];
assign
s_logisimBus42[16]
=
s_logisimBus88[16];
assign
s_logisimBus42[17]
=
s_logisimBus88[17];
assign
s_logisimBus42[18]
=
s_logisimBus88[18];
assign
s_logisimBus42[19]
=
s_logisimBus88[19];
assign
s_logisimBus42[20]
=
s_logisimBus88[20];
assign
s_logisimBus42[21]
=
s_logisimBus88[21];
assign
s_logisimBus42[22]
=
s_logisimBus88[22];
assign
s_logisimBus42[23]
=
s_logisimBus88[23];
assign
s_logisimBus42[24]
=
s_logisimBus88[24];
assign
s_logisimBus42[25]
=
s_logisimBus88[25];
assign
s_logisimBus42[26]
=
s_logisimBus88[26];
assign
s_logisimBus42[27]
=
s_logisimBus88[27];
assign
s_logisimBus42[28]
=
s_logisimBus88[28];
assign
s_logisimBus42[29]
=
s_logisimBus88[29];
assign
s_logisimBus42[30]
=
s_logisimBus88[30];
assign
s_logisimBus42[31]
=
s_logisimBus88[31];
assign
s_logisimBus42[32]
=
s_logisimBus88[31];
assign
s_logisimBus42[33]
=
s_logisimBus88[31];
assign
s_logisimBus42[34]
=
s_logisimBus88[31];
assign
s_logisimBus42[35]
=
s_logisimBus88[31];
assign
s_logisimBus42[36]
=
s_logisimBus88[31];
assign
s_logisimBus42[37]
=
s_logisimBus88[31];
assign
s_logisimBus42[38]
=
s_logisimBus88[31];
assign
s_logisimBus42[39]
=
s_logisimBus88[31];
assign
s_logisimBus42[40]
=
s_logisimBus88[31];
assign
s_logisimBus42[41]
=
s_logisimBus88[31];
assign
s_logisimBus42[42]
=
s_logisimBus88[31];
assign
s_logisimBus42[43]
=
s_logisimBus88[31];
assign
s_logisimBus42[44]
=
s_logisimBus88[31];
assign
s_logisimBus42[45]
=
s_logisimBus88[31];
assign
s_logisimBus42[46]
=
s_logisimBus88[31];
assign
s_logisimBus42[47]
=
s_logisimBus88[31];
assign
s_logisimBus42[48]
=
s_logisimBus88[31];
assign
s_logisimBus42[49]
=
s_logisimBus88[31];
assign
s_logisimBus42[50]
=
s_logisimBus88[31];
assign
s_logisimBus42[51]
=
s_logisimBus88[31];
assign
s_logisimBus42[52]
=
s_logisimBus88[31];
assign
s_logisimBus42[53]
=
s_logisimBus88[31];
assign
s_logisimBus42[54]
=
s_logisimBus88[31];
assign
s_logisimBus42[55]
=
s_logisimBus88[31];
assign
s_logisimBus42[56]
=
s_logisimBus88[31];
assign
s_logisimBus42[57]
=
s_logisimBus88[31];
assign
s_logisimBus42[58]
=
s_logisimBus88[31];
assign
s_logisimBus42[59]
=
s_logisimBus88[31];
assign
s_logisimBus42[60]
=
s_logisimBus88[31];
assign
s_logisimBus42[61]
=
s_logisimBus88[31];
assign
s_logisimBus42[62]
=
s_logisimBus88[31];
assign
s_logisimBus42[63]
=
s_logisimBus88[31];
assign
s_logisimNet2
=
~s_logisimNet44;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
AND_GATE_3_INPUTS
#(.BubblesMask(3'b000))
GATES_1
(.input1(s_logisimNet15),
.input2(1'b1),
.input3(s_logisimNet49),
.result(s_logisimNet71));
AND_GATE_3_INPUTS
#(.BubblesMask(3'b000))
GATES_2
(.input1(s_logisimNet54),
.input2(1'b1),
.input3(s_logisimNet86),
.result(s_logisimNet18));
OR_GATE
#(.BubblesMask(2'b00))
GATES_3
(.input1(s_logisimNet94),
.input2(s_logisimNet92),
.result(s_logisimNet33));
AND_GATE
#(.BubblesMask(2'b00))
GATES_4
(.input1(s_logisimNet2),
.input2(s_logisimNet97),
.result(s_logisimNet23));
AND_GATE
#(.BubblesMask(2'b00))
GATES_5
(.input1(s_logisimNet44),
.input2(s_logisimNet27),
.result(s_logisimNet73));
AND_GATE
#(.BubblesMask(2'b00))
GATES_6
(.input1(s_logisimNet94),
.input2(s_logisimNet14),
.result(s_logisimNet97));
AND_GATE
#(.BubblesMask(2'b00))
GATES_7
(.input1(s_logisimNet51),
.input2(s_logisimNet87),
.result(s_logisimNet15));
AND_GATE
#(.BubblesMask(2'b00))
GATES_8
(.input1(s_logisimNet20),
.input2(s_logisimNet91),
.result(s_logisimNet93));
AND_GATE
#(.BubblesMask(2'b00))
GATES_9
(.input1(s_logisimNet94),
.input2(s_logisimNet21),
.result(s_logisimNet82));
Multiplexer_bus_2
#(.nrOfBits(9))
PLEXERS_10
(.enable(1'b1),
.muxIn_0(s_logisimBus53[8:0]),
.muxIn_1(s_logisimBus24[8:0]),
.muxOut(s_logisimBus10[8:0]),
.sel(s_logisimNet92));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_11
(.enable(1'b1),
.muxIn_0(s_logisimBus61[31:0]),
.muxIn_1(s_logisimBus1[31:0]),
.muxOut(s_logisimBus65[31:0]),
.sel(s_logisimNet62));
Multiplexer_bus_2
#(.nrOfBits(5))
PLEXERS_12
(.enable(1'b1),
.muxIn_0(s_logisimBus9[15:11]),
.muxIn_1(s_logisimBus9[20:16]),
.muxOut(s_logisimBus37[4:0]),
.sel(s_logisimNet96));
Multiplexer_bus_2
#(.nrOfBits(5))
PLEXERS_13
(.enable(1'b1),
.muxIn_0(s_logisimBus37[4:0]),
.muxIn_1(s_logisimBus75[4:0]),
.muxOut(s_logisimBus6[4:0]),
.sel(s_logisimNet81));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_14
(.enable(1'b1),
.muxIn_0(s_logisimBus88[31:0]),
.muxIn_1(s_logisimBus38[31:0]),
.muxOut(s_logisimBus61[31:0]),
.sel(s_logisimNet58));
Multiplexer_bus_2
#(.nrOfBits(5))
PLEXERS_15
(.enable(1'b1),
.muxIn_0(s_logisimBus64[4:0]),
.muxIn_1(s_logisimBus6[4:0]),
.muxOut(s_logisimBus78[4:0]),
.sel(s_logisimNet91));
Multiplexer_bus_2
#(.nrOfBits(9))
PLEXERS_16
(.enable(1'b1),
.muxIn_0(s_logisimBus13[8:0]),
.muxIn_1(s_logisimBus30[8:0]),
.muxOut(s_logisimBus29[8:0]),
.sel(s_logisimNet23));
Multiplexer_bus_2
#(.nrOfBits(9))
PLEXERS_17
(.enable(1'b1),
.muxIn_0(s_logisimBus29[8:0]),
.muxIn_1(s_logisimBus30[8:0]),
.muxOut(s_logisimBus47[8:0]),
.sel(s_logisimNet73));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_18
(.enable(1'b1),
.muxIn_0(s_logisimBus12[31:0]),
.muxIn_1(s_logisimBus34[31:0]),
.muxOut(s_logisimBus11[31:0]),
.sel(s_logisimNet22));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_19
(.enable(1'b1),
.muxIn_0(s_logisimBus70[31:0]),
.muxIn_1(s_logisimBus4[31:0]),
.muxOut(s_logisimBus76[31:0]),
.sel(s_logisimNet81));
Multiplexer_bus_2
#(.nrOfBits(9))
PLEXERS_20
(.enable(1'b1),
.muxIn_0(s_logisimBus47[8:0]),
.muxIn_1(s_logisimBus9[8:0]),
.muxOut(s_logisimBus31[8:0]),
.sel(s_logisimNet82));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_21
(.enable(1'b1),
.muxIn_0(s_logisimBus11[31:0]),
.muxIn_1(s_logisimBus8[31:0]),
.muxOut(s_logisimBus56[31:0]),
.sel(s_logisimNet48));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_22
(.enable(1'b1),
.muxIn_0(s_logisimBus74[31:0]),
.muxIn_1(s_logisimBus3[31:0]),
.muxOut(s_logisimBus0[31:0]),
.sel(s_logisimNet48));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_23
(.enable(1'b1),
.muxIn_0(s_logisimBus65[31:0]),
.muxIn_1(s_logisimBus16[31:0]),
.muxOut(s_logisimBus70[31:0]),
.sel(s_logisimNet46));
Multiplexer_bus_2
#(.nrOfBits(9))
PLEXERS_24
(.enable(1'b1),
.muxIn_0(s_logisimBus13[8:0]),
.muxIn_1(s_logisimBus31[8:0]),
.muxOut(s_logisimBus67[8:0]),
.sel(s_logisimNet94));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_25
(.enable(1'b1),
.muxIn_0(s_logisimBus66[31:0]),
.muxIn_1(s_logisimBus69[31:0]),
.muxOut(s_logisimBus16[31:0]),
.sel(s_logisimNet84));
Multiplexer_bus_2
#(.nrOfBits(9))
PLEXERS_26
(.enable(1'b1),
.muxIn_0(s_logisimBus67[8:0]),
.muxIn_1(s_logisimBus74[8:0]),
.muxOut(s_logisimBus53[8:0]),
.sel(s_logisimNet89));
Adder
#(.extendedBits(10),
.nrOfBits(9))
ARITH_27
(.carryIn(1'b0),
.carryOut(),
.dataA(s_logisimBus13[8:0]),
.dataB(s_logisimBus79[8:0]),
.result(s_logisimBus24[8:0]));
Comparator
#(.nrOfBits(32),
.twosComplement(0))
ARITH_28
(.aEqualsB(s_logisimNet44),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus88[31:0]),
.dataB(s_logisimBus32[31:0]));
Adder
#(.extendedBits(10),
.nrOfBits(9))
ARITH_29
(.carryIn(1'b0),
.carryOut(),
.dataA(s_logisimBus13[8:0]),
.dataB(s_logisimBus9[8:0]),
.result(s_logisimBus30[8:0]));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
ALU_High
(.clock(s_logisimNet95),
.clockEnable(s_logisimNet94),
.d(s_logisimBus52[31:0]),
.q(s_logisimBus59[31:0]),
.reset(1'b0),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
ALU_Low
(.clock(s_logisimNet95),
.clockEnable(s_logisimNet94),
.d(s_logisimBus55[31:0]),
.q(s_logisimBus88[31:0]),
.reset(1'b0),
.tick(1'b1));
D_FLIPFLOP
#(.invertClockEnable(0))
MEMORY_32
(.clock(s_logisimNet95),
.d(s_logisimNet91),
.preset(1'b0),
.q(s_logisimNet54),
.qBar(),
.reset(1'b0),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(9))
MEMORY_33
(.clock(s_logisimNet95),
.clockEnable(s_logisimNet98),
.d(s_logisimBus13[8:0]),
.q(s_logisimBus17[8:0]),
.reset(1'b0),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
lo
(.clock(s_logisimNet95),
.clockEnable(s_logisimNet18),
.d(s_logisimBus88[31:0]),
.q(s_logisimBus69[31:0]),
.reset(s_logisimNet80),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
HI
(.clock(s_logisimNet95),
.clockEnable(s_logisimNet18),
.d(s_logisimBus59[31:0]),
.q(s_logisimBus66[31:0]),
.reset(s_logisimNet80),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
MEMORY_36
(.clock(s_logisimNet95),
.clockEnable(s_logisimNet87),
.d(s_logisimBus50[31:0]),
.q(s_logisimBus38[31:0]),
.reset(1'b0),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(9))
PC2
(.clock(s_logisimNet95),
.clockEnable(s_logisimNet33),
.d(s_logisimBus10[8:0]),
.q(s_logisimBus13[8:0]),
.reset(s_logisimNet80),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
data_read1
(.clock(s_logisimNet95),
.clockEnable(s_logisimNet98),
.d(s_logisimBus26[31:0]),
.q(s_logisimBus74[31:0]),
.reset(1'b0),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
IR
(.clock(s_logisimNet95),
.clockEnable(s_logisimNet92),
.d(s_logisimBus28[31:0]),
.q(s_logisimBus9[31:0]),
.reset(s_logisimNet80),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
data_read2
(.clock(s_logisimNet95),
.clockEnable(s_logisimNet98),
.d(s_logisimBus12[31:0]),
.q(s_logisimBus3[31:0]),
.reset(1'b0),
.tick(1'b1));
/*******************************************************************************
**
Here
all
sub-circuits
are
defined
**
*******************************************************************************/
right_shifter_2
right_shift
(.a(s_logisimBus42[63:0]),
.a_2_right_shift(s_logisimBus57[63:0]));
ALU
mainALU
(.a(s_logisimBus0[31:0]),
.aluop(s_logisimBus90[3:0]),
.b(s_logisimBus56[31:0]),
.clk(s_logisimNet95),
.done(s_logisimNet49),
.output_inc(s_logisimNet19),
.output_inverted(s_logisimNet19),
.res_high(s_logisimBus52[31:0]),
.res_low(s_logisimBus55[31:0]),
.rst(s_logisimNet80));
regfile
reg_file
(.Aread0(s_logisimBus9[25:21]),
.Aread1(s_logisimBus9[20:16]),
.Awrite(s_logisimBus78[4:0]),
.Dread0(s_logisimBus26[31:0]),
.Dread1(s_logisimBus12[31:0]),
.Dwrite(s_logisimBus76[31:0]),
.R1(s_logisimBus99[31:0]),
.R10(s_logisimBus108[31:0]),
.R11(s_logisimBus109[31:0]),
.R12(s_logisimBus110[31:0]),
.R13(s_logisimBus111[31:0]),
.R14(s_logisimBus112[31:0]),
.R15(s_logisimBus113[31:0]),
.R16(s_logisimBus114[31:0]),
.R17(s_logisimBus115[31:0]),
.R18(s_logisimBus116[31:0]),
.R19(s_logisimBus117[31:0]),
.R2(s_logisimBus100[31:0]),
.R20(s_logisimBus118[31:0]),
.R21(s_logisimBus119[31:0]),
.R22(s_logisimBus120[31:0]),
.R23(s_logisimBus121[31:0]),
.R24(s_logisimBus122[31:0]),
.R25(s_logisimBus123[31:0]),
.R26(s_logisimBus124[31:0]),
.R27(s_logisimBus125[31:0]),
.R28(s_logisimBus126[31:0]),
.R29(s_logisimBus127[31:0]),
.R3(s_logisimBus101[31:0]),
.R30(s_logisimBus128[31:0]),
.R31(s_logisimBus129[31:0]),
.R4(s_logisimBus102[31:0]),
.R5(s_logisimBus103[31:0]),
.R6(s_logisimBus104[31:0]),
.R7(s_logisimBus105[31:0]),
.R8(s_logisimBus106[31:0]),
.R9(s_logisimBus107[31:0]),
.clk(s_logisimNet95),
.rst(s_logisimNet80));
jtag_ram512
D_MEM
(.Addr(s_logisimBus57[8:0]),
.Din(s_logisimBus12[31:0]),
.Dout(s_logisimBus50[31:0]),
.Jen(s_logisimNet35),
.Jin(s_logisimBus39[31:0]),
.Jout(s_logisimBus83[31:0]),
.Wen(s_logisimNet71),
.clk(s_logisimNet95));
handle_inst_done
handle_done
(.aluop(s_logisimBus90[3:0]),
.clk(s_logisimNet95),
.done(s_logisimNet49),
.inst_done(s_logisimNet68),
.is_div(s_logisimNet86),
.is_mul(s_logisimNet40),
.rst(s_logisimNet80));
Control_Unit
controller
(.Opcode(s_logisimBus9[31:26]),
.aluop(s_logisimBus90[3:0]),
.beq(s_logisimNet27),
.bne(s_logisimNet14),
.funct(s_logisimBus9[5:0]),
.is_div(s_logisimNet86),
.is_jal(s_logisimNet81),
.is_jr(s_logisimNet89),
.is_mul(s_logisimNet40),
.jump(s_logisimNet21),
.lo_or_hi(s_logisimNet84),
.mem_to_reg(s_logisimNet58),
.mem_write(s_logisimNet51),
.mf(s_logisimNet46),
.reg_write(s_logisimNet20),
.regdst(s_logisimNet96),
.sll_control(s_logisimNet48),
.slti(s_logisimNet62),
.source_2(s_logisimNet22));
jtag_ram512
I_MEM
(.Addr(s_logisimBus13[8:0]),
.Din(32'd0),
.Dout(s_logisimBus28[31:0]),
.Jen(s_logisimNet35),
.Jin(s_logisimBus41[31:0]),
.Jout(s_logisimBus39[31:0]),
.Wen(1'b0),
.clk(s_logisimNet95));
Onehot
OneHT
(.Exec(s_logisimNet94),
.IDecode(s_logisimNet98),
.IFetch(s_logisimNet92),
.Instdone(s_logisimNet68),
.Mem(s_logisimNet87),
.WB(s_logisimNet91),
.clk(s_logisimNet95),
.rst(s_logisimNet80));
endmodule