/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
main
**
**
**
*****************************************************************************/
module
main(
Jen,
Jin,
Jout,
R1,
R10,
R11,
R12,
R13,
R14,
R15,
R16,
R17,
R18,
R19,
R2,
R20,
R21,
R22,
R23,
R24,
R25,
R26,
R27,
R28,
R29,
R3,
R30,
R31,
R4,
R5,
R6,
R7,
R8,
R9,
clk,
rst
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
Jen;
input
[31:0]
Jin;
input
clk;
input
rst;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
[31:0]
Jout;
output
[31:0]
R1;
output
[31:0]
R10;
output
[31:0]
R11;
output
[31:0]
R12;
output
[31:0]
R13;
output
[31:0]
R14;
output
[31:0]
R15;
output
[31:0]
R16;
output
[31:0]
R17;
output
[31:0]
R18;
output
[31:0]
R19;
output
[31:0]
R2;
output
[31:0]
R20;
output
[31:0]
R21;
output
[31:0]
R22;
output
[31:0]
R23;
output
[31:0]
R24;
output
[31:0]
R25;
output
[31:0]
R26;
output
[31:0]
R27;
output
[31:0]
R28;
output
[31:0]
R29;
output
[31:0]
R3;
output
[31:0]
R30;
output
[31:0]
R31;
output
[31:0]
R4;
output
[31:0]
R5;
output
[31:0]
R6;
output
[31:0]
R7;
output
[31:0]
R8;
output
[31:0]
R9;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[31:0]
s_logisimBus0;
wire
[31:0]
s_logisimBus1;
wire
[31:0]
s_logisimBus10;
wire
[31:0]
s_logisimBus15;
wire
[8:0]
s_logisimBus19;
wire
[31:0]
s_logisimBus2;
wire
[31:0]
s_logisimBus20;
wire
[4:0]
s_logisimBus21;
wire
[8:0]
s_logisimBus23;
wire
[31:0]
s_logisimBus24;
wire
[31:0]
s_logisimBus25;
wire
[31:0]
s_logisimBus26;
wire
[31:0]
s_logisimBus27;
wire
[31:0]
s_logisimBus28;
wire
[31:0]
s_logisimBus29;
wire
[31:0]
s_logisimBus3;
wire
[31:0]
s_logisimBus30;
wire
[31:0]
s_logisimBus31;
wire
[31:0]
s_logisimBus32;
wire
[31:0]
s_logisimBus33;
wire
[31:0]
s_logisimBus34;
wire
[31:0]
s_logisimBus35;
wire
[31:0]
s_logisimBus36;
wire
[31:0]
s_logisimBus37;
wire
[31:0]
s_logisimBus38;
wire
[31:0]
s_logisimBus39;
wire
[31:0]
s_logisimBus4;
wire
[31:0]
s_logisimBus40;
wire
[31:0]
s_logisimBus41;
wire
[31:0]
s_logisimBus42;
wire
[31:0]
s_logisimBus43;
wire
[31:0]
s_logisimBus44;
wire
[31:0]
s_logisimBus45;
wire
[31:0]
s_logisimBus46;
wire
[31:0]
s_logisimBus47;
wire
[31:0]
s_logisimBus48;
wire
[31:0]
s_logisimBus49;
wire
[8:0]
s_logisimBus5;
wire
[31:0]
s_logisimBus50;
wire
[31:0]
s_logisimBus51;
wire
[31:0]
s_logisimBus52;
wire
[31:0]
s_logisimBus53;
wire
[31:0]
s_logisimBus54;
wire
[31:0]
s_logisimBus55;
wire
[3:0]
s_logisimBus7;
wire
s_logisimNet11;
wire
s_logisimNet12;
wire
s_logisimNet17;
wire
s_logisimNet6;
wire
s_logisimNet9;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus3[31:0]
=
Jin;
assign
s_logisimNet12
=
Jen;
assign
s_logisimNet17
=
rst;
assign
s_logisimNet9
=
clk;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
Jout
=
s_logisimBus4[31:0];
assign
R1
=
s_logisimBus25[31:0];
assign
R10
=
s_logisimBus34[31:0];
assign
R11
=
s_logisimBus35[31:0];
assign
R12
=
s_logisimBus36[31:0];
assign
R13
=
s_logisimBus37[31:0];
assign
R14
=
s_logisimBus38[31:0];
assign
R15
=
s_logisimBus39[31:0];
assign
R16
=
s_logisimBus40[31:0];
assign
R17
=
s_logisimBus41[31:0];
assign
R18
=
s_logisimBus42[31:0];
assign
R19
=
s_logisimBus43[31:0];
assign
R2
=
s_logisimBus26[31:0];
assign
R20
=
s_logisimBus44[31:0];
assign
R21
=
s_logisimBus45[31:0];
assign
R22
=
s_logisimBus46[31:0];
assign
R23
=
s_logisimBus47[31:0];
assign
R24
=
s_logisimBus48[31:0];
assign
R25
=
s_logisimBus49[31:0];
assign
R26
=
s_logisimBus50[31:0];
assign
R27
=
s_logisimBus51[31:0];
assign
R28
=
s_logisimBus52[31:0];
assign
R29
=
s_logisimBus53[31:0];
assign
R3
=
s_logisimBus27[31:0];
assign
R30
=
s_logisimBus54[31:0];
assign
R31
=
s_logisimBus55[31:0];
assign
R4
=
s_logisimBus28[31:0];
assign
R5
=
s_logisimBus29[31:0];
assign
R6
=
s_logisimBus30[31:0];
assign
R7
=
s_logisimBus31[31:0];
assign
R8
=
s_logisimBus32[31:0];
assign
R9
=
s_logisimBus33[31:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus19[8:0]
=
{1'b0,
8'h01};
assign
s_logisimBus20[0]
=
s_logisimBus10[0];
assign
s_logisimBus20[1]
=
s_logisimBus10[1];
assign
s_logisimBus20[2]
=
s_logisimBus10[2];
assign
s_logisimBus20[3]
=
s_logisimBus10[3];
assign
s_logisimBus20[4]
=
s_logisimBus10[4];
assign
s_logisimBus20[5]
=
s_logisimBus10[5];
assign
s_logisimBus20[6]
=
s_logisimBus10[6];
assign
s_logisimBus20[7]
=
s_logisimBus10[7];
assign
s_logisimBus20[8]
=
s_logisimBus10[8];
assign
s_logisimBus20[9]
=
s_logisimBus10[9];
assign
s_logisimBus20[10]
=
s_logisimBus10[10];
assign
s_logisimBus20[11]
=
s_logisimBus10[11];
assign
s_logisimBus20[12]
=
s_logisimBus10[12];
assign
s_logisimBus20[13]
=
s_logisimBus10[13];
assign
s_logisimBus20[14]
=
s_logisimBus10[14];
assign
s_logisimBus20[15]
=
s_logisimBus10[15];
assign
s_logisimBus20[16]
=
s_logisimBus10[15];
assign
s_logisimBus20[17]
=
s_logisimBus10[15];
assign
s_logisimBus20[18]
=
s_logisimBus10[15];
assign
s_logisimBus20[19]
=
s_logisimBus10[15];
assign
s_logisimBus20[20]
=
s_logisimBus10[15];
assign
s_logisimBus20[21]
=
s_logisimBus10[15];
assign
s_logisimBus20[22]
=
s_logisimBus10[15];
assign
s_logisimBus20[23]
=
s_logisimBus10[15];
assign
s_logisimBus20[24]
=
s_logisimBus10[15];
assign
s_logisimBus20[25]
=
s_logisimBus10[15];
assign
s_logisimBus20[26]
=
s_logisimBus10[15];
assign
s_logisimBus20[27]
=
s_logisimBus10[15];
assign
s_logisimBus20[28]
=
s_logisimBus10[15];
assign
s_logisimBus20[29]
=
s_logisimBus10[15];
assign
s_logisimBus20[30]
=
s_logisimBus10[15];
assign
s_logisimBus20[31]
=
s_logisimBus10[15];
assign
s_logisimNet11
=
1'b0;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
Multiplexer_bus_2
#(.nrOfBits(5))
PLEXERS_1
(.enable(1'b1),
.muxIn_0(s_logisimBus10[15:11]),
.muxIn_1(s_logisimBus10[20:16]),
.muxOut(s_logisimBus21[4:0]),
.sel(s_logisimBus10[29]));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_2
(.enable(1'b1),
.muxIn_0(s_logisimBus1[31:0]),
.muxIn_1(s_logisimBus20[31:0]),
.muxOut(s_logisimBus24[31:0]),
.sel(s_logisimBus10[29]));
Adder
#(.extendedBits(10),
.nrOfBits(9))
ARITH_3
(.carryIn(1'b0),
.carryOut(),
.dataA(s_logisimBus19[8:0]),
.dataB(s_logisimBus5[8:0]),
.result(s_logisimBus23[8:0]));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(9))
PC
(.clock(s_logisimNet9),
.clockEnable(1'b1),
.d(s_logisimBus23[8:0]),
.q(s_logisimBus5[8:0]),
.reset(s_logisimNet17),
.tick(1'b1));
/*******************************************************************************
**
Here
all
sub-circuits
are
defined
**
*******************************************************************************/
ALU
mainALU
(.a(s_logisimBus0[31:0]),
.aluop(s_logisimBus7[3:0]),
.b(s_logisimBus24[31:0]),
.clk(s_logisimNet9),
.done(),
.output_inc(s_logisimNet11),
.output_inverted(s_logisimNet11),
.res_high(),
.res_low(s_logisimBus2[31:0]),
.rst(s_logisimNet17));
regfile
reg_file
(.Aread0(s_logisimBus10[25:21]),
.Aread1(s_logisimBus10[20:16]),
.Awrite(s_logisimBus21[4:0]),
.Dread0(s_logisimBus0[31:0]),
.Dread1(s_logisimBus1[31:0]),
.Dwrite(s_logisimBus2[31:0]),
.R1(s_logisimBus25[31:0]),
.R10(s_logisimBus34[31:0]),
.R11(s_logisimBus35[31:0]),
.R12(s_logisimBus36[31:0]),
.R13(s_logisimBus37[31:0]),
.R14(s_logisimBus38[31:0]),
.R15(s_logisimBus39[31:0]),
.R16(s_logisimBus40[31:0]),
.R17(s_logisimBus41[31:0]),
.R18(s_logisimBus42[31:0]),
.R19(s_logisimBus43[31:0]),
.R2(s_logisimBus26[31:0]),
.R20(s_logisimBus44[31:0]),
.R21(s_logisimBus45[31:0]),
.R22(s_logisimBus46[31:0]),
.R23(s_logisimBus47[31:0]),
.R24(s_logisimBus48[31:0]),
.R25(s_logisimBus49[31:0]),
.R26(s_logisimBus50[31:0]),
.R27(s_logisimBus51[31:0]),
.R28(s_logisimBus52[31:0]),
.R29(s_logisimBus53[31:0]),
.R3(s_logisimBus27[31:0]),
.R30(s_logisimBus54[31:0]),
.R31(s_logisimBus55[31:0]),
.R4(s_logisimBus28[31:0]),
.R5(s_logisimBus29[31:0]),
.R6(s_logisimBus30[31:0]),
.R7(s_logisimBus31[31:0]),
.R8(s_logisimBus32[31:0]),
.R9(s_logisimBus33[31:0]),
.clk(s_logisimNet9),
.rst(s_logisimNet17));
jtag_ram512
D_MEM
(.Addr(9'd0),
.Din(32'd0),
.Dout(),
.Jen(s_logisimNet12),
.Jin(s_logisimBus15[31:0]),
.Jout(s_logisimBus4[31:0]),
.Wen(1'b0),
.clk(s_logisimNet9));
jtag_ram512
I_MEM
(.Addr(s_logisimBus5[8:0]),
.Din(32'd0),
.Dout(s_logisimBus10[31:0]),
.Jen(s_logisimNet12),
.Jin(s_logisimBus3[31:0]),
.Jout(s_logisimBus15[31:0]),
.Wen(1'b0),
.clk(s_logisimNet9));
Control_Unit
Control
(.Opcode(s_logisimBus10[31:26]),
.aluop(s_logisimBus7[3:0]),
.funct(s_logisimBus10[5:0]));
endmodule