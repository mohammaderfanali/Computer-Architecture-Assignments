/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
divison
**
**
**
*****************************************************************************/
module
divison(
clk,
dividend,
divisor,
done,
quotient,
remainder,
rst,
start
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
clk;
input
[31:0]
dividend;
input
[31:0]
divisor;
input
rst;
input
start;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
done;
output
[31:0]
quotient;
output
[31:0]
remainder;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[31:0]
s_logisimBus1;
wire
[31:0]
s_logisimBus13;
wire
[31:0]
s_logisimBus14;
wire
[6:0]
s_logisimBus15;
wire
[31:0]
s_logisimBus16;
wire
[31:0]
s_logisimBus17;
wire
[31:0]
s_logisimBus20;
wire
[31:0]
s_logisimBus22;
wire
[31:0]
s_logisimBus23;
wire
[6:0]
s_logisimBus24;
wire
[31:0]
s_logisimBus28;
wire
[31:0]
s_logisimBus29;
wire
[31:0]
s_logisimBus3;
wire
[31:0]
s_logisimBus30;
wire
[6:0]
s_logisimBus31;
wire
[31:0]
s_logisimBus4;
wire
[31:0]
s_logisimBus5;
wire
[6:0]
s_logisimBus6;
wire
[6:0]
s_logisimBus7;
wire
[31:0]
s_logisimBus8;
wire
s_logisimNet0;
wire
s_logisimNet10;
wire
s_logisimNet11;
wire
s_logisimNet12;
wire
s_logisimNet18;
wire
s_logisimNet19;
wire
s_logisimNet2;
wire
s_logisimNet21;
wire
s_logisimNet25;
wire
s_logisimNet26;
wire
s_logisimNet27;
wire
s_logisimNet9;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus13[31:0]
=
divisor;
assign
s_logisimBus17[31:0]
=
dividend;
assign
s_logisimNet11
=
start;
assign
s_logisimNet18
=
clk;
assign
s_logisimNet21
=
rst;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
done
=
s_logisimNet12;
assign
quotient
=
s_logisimBus5[31:0];
assign
remainder
=
s_logisimBus3[31:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus6[6:0]
=
{3'b000,
4'h0};
assign
s_logisimBus7[6:0]
=
{3'b010,
4'h0};
assign
s_logisimBus8[31:0]
=
32'h00000001;
assign
s_logisimNet19
=
1'b0;
assign
s_logisimBus16[31:0]
=
32'h00000000;
assign
s_logisimBus31[6:0]
=
{3'b000,
4'h0};
assign
s_logisimNet25
=
~s_logisimNet2;
assign
s_logisimNet9
=
~s_logisimNet10;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
OR_GATE_BUS
#(.BubblesMask(2'b00),
.NrOfBits(32))
GATES_1
(.input1(s_logisimBus1[31:0]),
.input2(s_logisimBus8[31:0]),
.result(s_logisimBus23[31:0]));
OR_GATE
#(.BubblesMask(2'b00))
GATES_2
(.input1(s_logisimNet11),
.input2(s_logisimNet2),
.result(s_logisimNet26));
OR_GATE
#(.BubblesMask(2'b00))
GATES_3
(.input1(s_logisimNet11),
.input2(s_logisimNet25),
.result(s_logisimNet0));
OR_GATE
#(.BubblesMask(2'b00))
GATES_4
(.input1(s_logisimNet12),
.input2(s_logisimNet2),
.result(s_logisimNet27));
Multiplexer_bus_2
#(.nrOfBits(7))
PLEXERS_5
(.enable(1'b1),
.muxIn_0(s_logisimBus6[6:0]),
.muxIn_1(s_logisimBus7[6:0]),
.muxOut(s_logisimBus15[6:0]),
.sel(s_logisimNet11));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_6
(.enable(1'b1),
.muxIn_0(s_logisimBus20[31:0]),
.muxIn_1(s_logisimBus17[31:0]),
.muxOut(s_logisimBus30[31:0]),
.sel(s_logisimNet11));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_7
(.enable(1'b1),
.muxIn_0(s_logisimBus1[31:0]),
.muxIn_1(s_logisimBus23[31:0]),
.muxOut(s_logisimBus20[31:0]),
.sel(s_logisimNet9));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_8
(.enable(1'b1),
.muxIn_0(s_logisimBus4[31:0]),
.muxIn_1(s_logisimBus28[31:0]),
.muxOut(s_logisimBus22[31:0]),
.sel(s_logisimNet9));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_9
(.enable(1'b1),
.muxIn_0(s_logisimBus22[31:0]),
.muxIn_1(s_logisimBus16[31:0]),
.muxOut(s_logisimBus29[31:0]),
.sel(s_logisimNet11));
Subtractor
#(.extendedBits(33),
.nrOfBits(32))
ARITH_10
(.borrowIn(1'b0),
.borrowOut(),
.dataA(s_logisimBus4[31:0]),
.dataB(s_logisimBus14[31:0]),
.result(s_logisimBus28[31:0]));
Comparator
#(.nrOfBits(7),
.twosComplement(0))
ARITH_11
(.aEqualsB(s_logisimNet2),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus31[6:0]),
.dataB(s_logisimBus24[6:0]));
Comparator
#(.nrOfBits(32),
.twosComplement(0))
ARITH_12
(.aEqualsB(),
.aGreaterThanB(s_logisimNet10),
.aLessThanB(),
.dataA(s_logisimBus14[31:0]),
.dataB(s_logisimBus4[31:0]));
LogisimCounter
#(.invertClock(0),
.maxVal({3'b111,
4'hF}),
.mode(0),
.width(7))
MEMORY_13
(.clear(1'b0),
.clock(s_logisimNet18),
.compareOut(),
.countValue(s_logisimBus24[6:0]),
.enable(1'b1),
.load(s_logisimNet26),
.loadData(s_logisimBus15[6:0]),
.tick(1'b1),
.upNotDown(s_logisimNet19));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
q
(.clock(s_logisimNet18),
.clockEnable(s_logisimNet0),
.d(s_logisimBus30[31:0]),
.q(s_logisimBus5[31:0]),
.reset(s_logisimNet21),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
a
(.clock(s_logisimNet18),
.clockEnable(s_logisimNet0),
.d(s_logisimBus29[31:0]),
.q(s_logisimBus3[31:0]),
.reset(s_logisimNet21),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
b
(.clock(s_logisimNet18),
.clockEnable(s_logisimNet11),
.d(s_logisimBus13[31:0]),
.q(s_logisimBus14[31:0]),
.reset(s_logisimNet21),
.tick(1'b1));
D_FLIPFLOP
#(.invertClockEnable(0))
MEMORY_17
(.clock(s_logisimNet18),
.d(s_logisimNet27),
.preset(1'b0),
.q(s_logisimNet12),
.qBar(),
.reset(s_logisimNet11),
.tick(1'b1));
/*******************************************************************************
**
Here
all
sub-circuits
are
defined
**
*******************************************************************************/
shift
shift_1
(.a(s_logisimBus3[31:0]),
.new_a(s_logisimBus4[31:0]),
.new_q(s_logisimBus1[31:0]),
.q(s_logisimBus5[31:0]));
endmodule