/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
Carry_Select_Adder
**
**
**
*****************************************************************************/
module
Carry_Select_Adder(
Carry_in,
Carry_out,
Sum,
a,
b
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
Carry_in;
input
[31:0]
a;
input
[31:0]
b;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
Carry_out;
output
[31:0]
Sum;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[7:0]
s_logisimBus11;
wire
[7:0]
s_logisimBus16;
wire
[7:0]
s_logisimBus2;
wire
[7:0]
s_logisimBus21;
wire
[7:0]
s_logisimBus30;
wire
[7:0]
s_logisimBus31;
wire
[31:0]
s_logisimBus35;
wire
[31:0]
s_logisimBus4;
wire
[31:0]
s_logisimBus9;
wire
s_logisimNet0;
wire
s_logisimNet13;
wire
s_logisimNet14;
wire
s_logisimNet15;
wire
s_logisimNet17;
wire
s_logisimNet20;
wire
s_logisimNet22;
wire
s_logisimNet24;
wire
s_logisimNet29;
wire
s_logisimNet32;
wire
s_logisimNet33;
wire
s_logisimNet34;
wire
s_logisimNet36;
wire
s_logisimNet37;
wire
s_logisimNet5;
wire
s_logisimNet6;
wire
s_logisimNet8;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus35[31:0]
=
a;
assign
s_logisimBus4[31:0]
=
b;
assign
s_logisimNet20
=
Carry_in;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
Carry_out
=
s_logisimNet34;
assign
Sum
=
s_logisimBus9[31:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimNet6
=
1'b0;
assign
s_logisimNet32
=
1'b0;
assign
s_logisimNet36
=
1'b0;
assign
s_logisimNet15
=
1'b1;
assign
s_logisimNet33
=
1'b1;
assign
s_logisimNet37
=
1'b1;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
Multiplexer_bus_2
#(.nrOfBits(8))
PLEXERS_1
(.enable(1'b1),
.muxIn_0(s_logisimBus11[7:0]),
.muxIn_1(s_logisimBus21[7:0]),
.muxOut(s_logisimBus9[31:24]),
.sel(s_logisimNet24));
Multiplexer_bus_2
#(.nrOfBits(8))
PLEXERS_2
(.enable(1'b1),
.muxIn_0(s_logisimBus31[7:0]),
.muxIn_1(s_logisimBus30[7:0]),
.muxOut(s_logisimBus9[23:16]),
.sel(s_logisimNet0));
Multiplexer_bus_2
#(.nrOfBits(8))
PLEXERS_3
(.enable(1'b1),
.muxIn_0(s_logisimBus2[7:0]),
.muxIn_1(s_logisimBus16[7:0]),
.muxOut(s_logisimBus9[15:8]),
.sel(s_logisimNet8));
Multiplexer_2
PLEXERS_4
(.enable(1'b1),
.muxIn_0(s_logisimNet5),
.muxIn_1(s_logisimNet29),
.muxOut(s_logisimNet34),
.sel(s_logisimNet24));
Multiplexer_2
PLEXERS_5
(.enable(1'b1),
.muxIn_0(s_logisimNet14),
.muxIn_1(s_logisimNet13),
.muxOut(s_logisimNet24),
.sel(s_logisimNet0));
Multiplexer_2
PLEXERS_6
(.enable(1'b1),
.muxIn_0(s_logisimNet22),
.muxIn_1(s_logisimNet17),
.muxOut(s_logisimNet0),
.sel(s_logisimNet8));
Adder
#(.extendedBits(9),
.nrOfBits(8))
ARITH_7
(.carryIn(s_logisimNet32),
.carryOut(s_logisimNet14),
.dataA(s_logisimBus35[23:16]),
.dataB(s_logisimBus4[23:16]),
.result(s_logisimBus31[7:0]));
Adder
#(.extendedBits(9),
.nrOfBits(8))
ARITH_8
(.carryIn(s_logisimNet36),
.carryOut(s_logisimNet22),
.dataA(s_logisimBus35[15:8]),
.dataB(s_logisimBus4[15:8]),
.result(s_logisimBus2[7:0]));
Adder
#(.extendedBits(9),
.nrOfBits(8))
ARITH_9
(.carryIn(s_logisimNet6),
.carryOut(s_logisimNet5),
.dataA(s_logisimBus35[31:24]),
.dataB(s_logisimBus4[31:24]),
.result(s_logisimBus11[7:0]));
Adder
#(.extendedBits(9),
.nrOfBits(8))
ARITH_10
(.carryIn(s_logisimNet20),
.carryOut(s_logisimNet8),
.dataA(s_logisimBus35[7:0]),
.dataB(s_logisimBus4[7:0]),
.result(s_logisimBus9[7:0]));
Adder
#(.extendedBits(9),
.nrOfBits(8))
ARITH_11
(.carryIn(s_logisimNet33),
.carryOut(s_logisimNet13),
.dataA(s_logisimBus35[23:16]),
.dataB(s_logisimBus4[23:16]),
.result(s_logisimBus30[7:0]));
Adder
#(.extendedBits(9),
.nrOfBits(8))
ARITH_12
(.carryIn(s_logisimNet37),
.carryOut(s_logisimNet17),
.dataA(s_logisimBus35[15:8]),
.dataB(s_logisimBus4[15:8]),
.result(s_logisimBus16[7:0]));
Adder
#(.extendedBits(9),
.nrOfBits(8))
ARITH_13
(.carryIn(s_logisimNet15),
.carryOut(s_logisimNet29),
.dataA(s_logisimBus35[31:24]),
.dataB(s_logisimBus4[31:24]),
.result(s_logisimBus21[7:0]));
endmodule