/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
multiply
**
**
**
*****************************************************************************/
module
multiply(
a,
b,
clk,
done,
res_high,
res_low,
rst,
start
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[31:0]
a;
input
[31:0]
b;
input
clk;
input
rst;
input
start;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
done;
output
[31:0]
res_high;
output
[31:0]
res_low;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[31:0]
s_logisimBus0;
wire
[31:0]
s_logisimBus12;
wire
[31:0]
s_logisimBus13;
wire
[31:0]
s_logisimBus14;
wire
[31:0]
s_logisimBus15;
wire
[63:0]
s_logisimBus16;
wire
[31:0]
s_logisimBus20;
wire
[31:0]
s_logisimBus23;
wire
[31:0]
s_logisimBus25;
wire
[31:0]
s_logisimBus26;
wire
[6:0]
s_logisimBus27;
wire
[63:0]
s_logisimBus31;
wire
[6:0]
s_logisimBus32;
wire
[63:0]
s_logisimBus33;
wire
[31:0]
s_logisimBus35;
wire
[6:0]
s_logisimBus36;
wire
[31:0]
s_logisimBus39;
wire
[31:0]
s_logisimBus40;
wire
[63:0]
s_logisimBus42;
wire
[6:0]
s_logisimBus43;
wire
[6:0]
s_logisimBus6;
wire
[31:0]
s_logisimBus8;
wire
[31:0]
s_logisimBus9;
wire
s_logisimNet1;
wire
s_logisimNet10;
wire
s_logisimNet17;
wire
s_logisimNet18;
wire
s_logisimNet2;
wire
s_logisimNet21;
wire
s_logisimNet22;
wire
s_logisimNet24;
wire
s_logisimNet28;
wire
s_logisimNet29;
wire
s_logisimNet3;
wire
s_logisimNet34;
wire
s_logisimNet38;
wire
s_logisimNet7;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus0[31:0]
=
a;
assign
s_logisimBus8[31:0]
=
b;
assign
s_logisimNet18
=
rst;
assign
s_logisimNet2
=
clk;
assign
s_logisimNet34
=
start;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
done
=
s_logisimNet7;
assign
res_high
=
s_logisimBus15[31:0];
assign
res_low
=
s_logisimBus31[31:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus25[29:0]
=
{2'b00,
28'h0000000};
assign
s_logisimBus12[31:0]
=
32'h00000000;
assign
s_logisimBus13[31:0]
=
32'h00000000;
assign
s_logisimBus6[6:0]
=
{3'b000,
4'h0};
assign
s_logisimBus36[6:0]
=
{3'b001,
4'h0};
assign
s_logisimNet17
=
1'b0;
assign
s_logisimBus43[6:0]
=
{3'b000,
4'h0};
assign
s_logisimBus42[63:32]
=
32'h00000000;
assign
s_logisimBus20[31:0]
=
32'h00000000;
assign
s_logisimBus31[63:32]
=
32'h00000000;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
OR_GATE_BUS
#(.BubblesMask(2'b00),
.NrOfBits(32))
GATES_1
(.input1(s_logisimBus16[31:0]),
.input2(s_logisimBus25[31:0]),
.result(s_logisimBus9[31:0]));
OR_GATE
#(.BubblesMask(2'b00))
GATES_2
(.input1(s_logisimNet34),
.input2(s_logisimNet1),
.result(s_logisimNet29));
OR_GATE
#(.BubblesMask(2'b00))
GATES_3
(.input1(s_logisimNet34),
.input2(s_logisimNet10),
.result(s_logisimNet28));
OR_GATE
#(.BubblesMask(2'b00))
GATES_4
(.input1(s_logisimNet7),
.input2(s_logisimNet1),
.result(s_logisimNet38));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_5
(.enable(1'b1),
.muxIn_0(s_logisimBus9[31:0]),
.muxIn_1(s_logisimBus12[31:0]),
.muxOut(s_logisimBus35[31:0]),
.sel(s_logisimNet34));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_6
(.enable(1'b1),
.muxIn_0(s_logisimBus23[31:0]),
.muxIn_1(s_logisimBus13[31:0]),
.muxOut(s_logisimBus26[31:0]),
.sel(s_logisimNet34));
Multiplexer_bus_2
#(.nrOfBits(7))
PLEXERS_7
(.enable(1'b1),
.muxIn_0(s_logisimBus6[6:0]),
.muxIn_1(s_logisimBus36[6:0]),
.muxOut(s_logisimBus32[6:0]),
.sel(s_logisimNet34));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_8
(.enable(1'b1),
.muxIn_0(s_logisimBus33[31:0]),
.muxIn_1(s_logisimBus8[31:0]),
.muxOut(s_logisimBus39[31:0]),
.sel(s_logisimNet34));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_9
(.enable(1'b1),
.muxIn_0(s_logisimBus20[31:0]),
.muxIn_1(s_logisimBus0[31:0]),
.muxOut(s_logisimBus14[31:0]),
.sel(s_logisimBus42[0]));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_10
(.enable(1'b1),
.muxIn_0(s_logisimBus20[31:0]),
.muxIn_1(s_logisimBus0[31:0]),
.muxOut(s_logisimBus40[31:0]),
.sel(s_logisimBus42[1]));
Comparator
#(.nrOfBits(7),
.twosComplement(0))
ARITH_11
(.aEqualsB(s_logisimNet1),
.aGreaterThanB(),
.aLessThanB(s_logisimNet10),
.dataA(s_logisimBus43[6:0]),
.dataB(s_logisimBus27[6:0]));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
MEMORY_12
(.clock(s_logisimNet2),
.clockEnable(s_logisimNet28),
.d(s_logisimBus35[31:0]),
.q(s_logisimBus31[31:0]),
.reset(s_logisimNet18),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
MEMORY_13
(.clock(s_logisimNet2),
.clockEnable(s_logisimNet28),
.d(s_logisimBus26[31:0]),
.q(s_logisimBus15[31:0]),
.reset(s_logisimNet18),
.tick(1'b1));
LogisimCounter
#(.invertClock(0),
.maxVal({3'b111,
4'hF}),
.mode(0),
.width(7))
MEMORY_14
(.clear(1'b0),
.clock(s_logisimNet2),
.compareOut(),
.countValue(s_logisimBus27[6:0]),
.enable(1'b1),
.load(s_logisimNet29),
.loadData(s_logisimBus32[6:0]),
.tick(1'b1),
.upNotDown(s_logisimNet17));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
MEMORY_15
(.clock(s_logisimNet2),
.clockEnable(s_logisimNet28),
.d(s_logisimBus39[31:0]),
.q(s_logisimBus42[31:0]),
.reset(s_logisimNet18),
.tick(1'b1));
D_FLIPFLOP
#(.invertClockEnable(0))
MEMORY_16
(.clock(s_logisimNet2),
.d(s_logisimNet38),
.preset(1'b0),
.q(s_logisimNet7),
.qBar(),
.reset(s_logisimNet34),
.tick(1'b1));
/*******************************************************************************
**
Here
all
sub-circuits
are
defined
**
*******************************************************************************/
right_shifter_2
right_shifter_2_2
(.a(s_logisimBus31[63:0]),
.a_2_right_shift(s_logisimBus16[63:0]));
Carry_Save_Adder
CSA
(.S0(s_logisimBus25[30]),
.S1(s_logisimBus25[31]),
.a(s_logisimBus15[31:0]),
.b(s_logisimBus14[31:0]),
.c(s_logisimBus40[31:0]),
.new_S(s_logisimBus23[31:0]));
right_shifter_2
right_shifter_2_1
(.a(s_logisimBus42[63:0]),
.a_2_right_shift(s_logisimBus33[63:0]));
endmodule