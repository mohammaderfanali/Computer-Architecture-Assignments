/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
handle_start
**
**
**
*****************************************************************************/
module
handle_start(
a,
aluop,
b,
clk,
rst,
start
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[31:0]
a;
input
[3:0]
aluop;
input
[31:0]
b;
input
clk;
input
rst;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
start;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[31:0]
s_logisimBus10;
wire
[3:0]
s_logisimBus16;
wire
[31:0]
s_logisimBus19;
wire
[31:0]
s_logisimBus2;
wire
[3:0]
s_logisimBus4;
wire
[31:0]
s_logisimBus5;
wire
[3:0]
s_logisimBus8;
wire
s_logisimNet0;
wire
s_logisimNet1;
wire
s_logisimNet11;
wire
s_logisimNet12;
wire
s_logisimNet13;
wire
s_logisimNet14;
wire
s_logisimNet15;
wire
s_logisimNet17;
wire
s_logisimNet18;
wire
s_logisimNet20;
wire
s_logisimNet3;
wire
s_logisimNet6;
wire
s_logisimNet7;
wire
s_logisimNet9;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus10[31:0]
=
b;
assign
s_logisimBus2[31:0]
=
a;
assign
s_logisimBus8[3:0]
=
aluop;
assign
s_logisimNet1
=
clk;
assign
s_logisimNet11
=
rst;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
start
=
s_logisimNet15;
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus4[3:0]
=
4'h2;
assign
s_logisimBus16[3:0]
=
4'h3;
assign
s_logisimNet7
=
1'b1;
assign
s_logisimNet20
=
1'b1;
assign
s_logisimNet14
=
~s_logisimNet9;
assign
s_logisimNet0
=
~s_logisimNet18;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
OR_GATE
#(.BubblesMask(2'b00))
GATES_1
(.input1(s_logisimNet14),
.input2(s_logisimNet0),
.result(s_logisimNet3));
AND_GATE
#(.BubblesMask(2'b00))
GATES_2
(.input1(s_logisimNet3),
.input2(s_logisimNet13),
.result(s_logisimNet6));
OR_GATE
#(.BubblesMask(2'b00))
GATES_3
(.input1(s_logisimNet17),
.input2(s_logisimNet12),
.result(s_logisimNet13));
Comparator
#(.nrOfBits(4),
.twosComplement(1))
ARITH_4
(.aEqualsB(s_logisimNet17),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus8[3:0]),
.dataB(s_logisimBus4[3:0]));
Comparator
#(.nrOfBits(4),
.twosComplement(1))
ARITH_5
(.aEqualsB(s_logisimNet12),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus8[3:0]),
.dataB(s_logisimBus16[3:0]));
Comparator
#(.nrOfBits(32),
.twosComplement(1))
ARITH_6
(.aEqualsB(s_logisimNet9),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus19[31:0]),
.dataB(s_logisimBus2[31:0]));
Comparator
#(.nrOfBits(32),
.twosComplement(1))
ARITH_7
(.aEqualsB(s_logisimNet18),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus5[31:0]),
.dataB(s_logisimBus10[31:0]));
D_FLIPFLOP
#(.invertClockEnable(0))
MEMORY_8
(.clock(s_logisimNet1),
.d(s_logisimNet6),
.preset(1'b0),
.q(s_logisimNet15),
.qBar(),
.reset(s_logisimNet11),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
MEMORY_9
(.clock(s_logisimNet1),
.clockEnable(s_logisimNet20),
.d(s_logisimBus2[31:0]),
.q(s_logisimBus19[31:0]),
.reset(s_logisimNet11),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
MEMORY_10
(.clock(s_logisimNet1),
.clockEnable(s_logisimNet7),
.d(s_logisimBus10[31:0]),
.q(s_logisimBus5[31:0]),
.reset(s_logisimNet11),
.tick(1'b1));
endmodule