/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
handle_inst_done
**
**
**
*****************************************************************************/
module
handle_inst_done(
aluop,
clk,
done,
inst_done,
is_div,
is_mul,
rst
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[3:0]
aluop;
input
clk;
input
done;
input
is_div;
input
is_mul;
input
rst;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
inst_done;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[3:0]
s_logisimBus11;
wire
[3:0]
s_logisimBus2;
wire
s_logisimNet0;
wire
s_logisimNet1;
wire
s_logisimNet10;
wire
s_logisimNet12;
wire
s_logisimNet13;
wire
s_logisimNet3;
wire
s_logisimNet4;
wire
s_logisimNet5;
wire
s_logisimNet6;
wire
s_logisimNet7;
wire
s_logisimNet8;
wire
s_logisimNet9;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus2[3:0]
=
aluop;
assign
s_logisimNet1
=
is_mul;
assign
s_logisimNet4
=
clk;
assign
s_logisimNet5
=
is_div;
assign
s_logisimNet7
=
rst;
assign
s_logisimNet9
=
done;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
inst_done
=
s_logisimNet10;
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimNet8
=
1'b0;
assign
s_logisimNet13
=
1'b1;
assign
s_logisimNet3
=
~s_logisimNet6;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
OR_GATE
#(.BubblesMask(2'b00))
GATES_1
(.input1(s_logisimNet1),
.input2(s_logisimNet5),
.result(s_logisimNet12));
AND_GATE
#(.BubblesMask(2'b00))
GATES_2
(.input1(s_logisimNet3),
.input2(s_logisimNet12),
.result(s_logisimNet0));
Multiplexer_2
PLEXERS_3
(.enable(1'b1),
.muxIn_0(s_logisimNet9),
.muxIn_1(s_logisimNet8),
.muxOut(s_logisimNet10),
.sel(s_logisimNet0));
Comparator
#(.nrOfBits(4),
.twosComplement(0))
ARITH_4
(.aEqualsB(s_logisimNet6),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus11[3:0]),
.dataB(s_logisimBus2[3:0]));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(4))
MEMORY_5
(.clock(s_logisimNet4),
.clockEnable(s_logisimNet13),
.d(s_logisimBus2[3:0]),
.q(s_logisimBus11[3:0]),
.reset(s_logisimNet7),
.tick(1'b1));
endmodule