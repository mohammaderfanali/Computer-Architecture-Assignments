/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
Control_Unit
**
**
**
*****************************************************************************/
module
Control_Unit(
Opcode,
aluop,
funct
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[5:0]
Opcode;
input
[5:0]
funct;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
[3:0]
aluop;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[3:0]
s_logisimBus13;
wire
[5:0]
s_logisimBus18;
wire
[5:0]
s_logisimBus20;
wire
[3:0]
s_logisimBus21;
wire
[3:0]
s_logisimBus5;
wire
s_logisimNet0;
wire
s_logisimNet1;
wire
s_logisimNet10;
wire
s_logisimNet11;
wire
s_logisimNet12;
wire
s_logisimNet14;
wire
s_logisimNet15;
wire
s_logisimNet16;
wire
s_logisimNet17;
wire
s_logisimNet19;
wire
s_logisimNet2;
wire
s_logisimNet22;
wire
s_logisimNet23;
wire
s_logisimNet24;
wire
s_logisimNet3;
wire
s_logisimNet4;
wire
s_logisimNet6;
wire
s_logisimNet7;
wire
s_logisimNet8;
wire
s_logisimNet9;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus18[5:0]
=
Opcode;
assign
s_logisimBus20[5:0]
=
funct;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
aluop
=
s_logisimBus13[3:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus21[3:0]
=
4'h0;
assign
s_logisimNet6
=
~s_logisimBus20[5];
assign
s_logisimNet7
=
~s_logisimBus20[5];
assign
s_logisimNet8
=
~s_logisimBus20[1];
assign
s_logisimNet22
=
~s_logisimBus20[0];
assign
s_logisimNet23
=
~s_logisimBus20[1];
assign
s_logisimNet24
=
~s_logisimBus20[2];
assign
s_logisimNet9
=
~s_logisimBus20[0];
assign
s_logisimBus5[3]
=
~s_logisimBus20[5];
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
AND_GATE
#(.BubblesMask(2'b00))
GATES_1
(.input1(s_logisimBus20[1]),
.input2(s_logisimBus20[2]),
.result(s_logisimBus5[1]));
AND_GATE
#(.BubblesMask(2'b00))
GATES_2
(.input1(s_logisimBus20[2]),
.input2(s_logisimBus20[5]),
.result(s_logisimBus5[2]));
AND_GATE_4_INPUTS
#(.BubblesMask(4'h0))
GATES_3
(.input1(s_logisimBus20[2]),
.input2(s_logisimNet6),
.input3(s_logisimBus20[1]),
.input4(s_logisimBus20[0]),
.result(s_logisimNet12));
AND_GATE_4_INPUTS
#(.BubblesMask(4'h0))
GATES_4
(.input1(s_logisimBus20[2]),
.input2(s_logisimNet7),
.input3(s_logisimNet8),
.input4(s_logisimNet22),
.result(s_logisimNet17));
AND_GATE_4_INPUTS
#(.BubblesMask(4'h0))
GATES_5
(.input1(s_logisimBus20[2]),
.input2(s_logisimBus20[5]),
.input3(s_logisimNet23),
.input4(s_logisimBus20[0]),
.result(s_logisimNet14));
AND_GATE_4_INPUTS
#(.BubblesMask(4'h0))
GATES_6
(.input1(s_logisimBus20[5]),
.input2(s_logisimNet24),
.input3(s_logisimBus20[1]),
.input4(s_logisimNet9),
.result(s_logisimNet19));
OR_GATE_4_INPUTS
#(.BubblesMask(4'h0))
GATES_7
(.input1(s_logisimNet12),
.input2(s_logisimNet17),
.input3(s_logisimNet14),
.input4(s_logisimNet19),
.result(s_logisimBus5[0]));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_8
(.enable(1'b1),
.muxIn_0(s_logisimBus5[3:0]),
.muxIn_1(s_logisimBus21[3:0]),
.muxOut(s_logisimBus13[3:0]),
.sel(s_logisimBus18[3]));
endmodule