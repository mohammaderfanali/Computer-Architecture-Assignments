/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
OR_GATE
**
**
**
*****************************************************************************/
module
OR_GATE(
input1,
input2,
result
);
/*******************************************************************************
**
Here
all
module
parameters
are
defined
with
a
dummy
value
**
*******************************************************************************/
parameter
[64:0]
BubblesMask
=
1;
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
input1;
input
input2;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
result;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
s_realInput1;
wire
s_realInput2;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
the
bubbles
are
processed
**
*******************************************************************************/
assign
s_realInput1
=
(BubblesMask[0]
==
1'b0)
?
input1
:
~input1;
assign
s_realInput2
=
(BubblesMask[1]
==
1'b0)
?
input2
:
~input2;
/*******************************************************************************
**
Here
the
functionality
is
defined
**
*******************************************************************************/
assign
result
=
s_realInput1|
s_realInput2;
endmodule