/******************************************************************************
 ** Logisim-evolution goes FPGA automatic generated Verilog code             **
 ** https://github.com/logisim-evolution/                                    **
 **                                                                          **
 ** Component : sign_extended                                                **
 **                                                                          **
 *****************************************************************************/

module sign_extended( a,
                      a_extend,
                      sign );

   /*******************************************************************************
   ** The inputs are defined here                                                **
   *******************************************************************************/
   input [31:0] a;
   input        sign;

   /*******************************************************************************
   ** The outputs are defined here                                               **
   *******************************************************************************/
   output [63:0] a_extend;

   /*******************************************************************************
   ** The wires are defined here                                                 **
   *******************************************************************************/
   wire [31:0] s_logisimBus1;
   wire [31:0] s_logisimBus4;
   wire [63:0] s_logisimBus6;
   wire [31:0] s_logisimBus7;
   wire [31:0] s_logisimBus8;
   wire        s_logisimNet3;
   wire        s_logisimNet5;

   /*******************************************************************************
   ** The module functionality is described here                                 **
   *******************************************************************************/

   /*******************************************************************************
   ** Here all input connections are defined                                     **
   *******************************************************************************/
   assign s_logisimBus6[31:0] = a;
   assign s_logisimNet5       = sign;

   /*******************************************************************************
   ** Here all output connections are defined                                    **
   *******************************************************************************/
   assign a_extend = s_logisimBus6[63:0];

   /*******************************************************************************
   ** Here all in-lined components are defined                                   **
   *******************************************************************************/

   // Constant
   assign  s_logisimBus4[31:0]  =  32'h00000000;


   // Constant
   assign  s_logisimBus7[31:0]  =  32'hFFFFFFFF;


   // Constant
   assign  s_logisimBus8[31:0]  =  32'h00000000;


   /*******************************************************************************
   ** Here all normal components are defined                                     **
   *******************************************************************************/
   Multiplexer_bus_2 #(.nrOfBits(32))
      PLEXERS_1 (.enable(1'b1),
                 .muxIn_0(s_logisimBus4[31:0]),
                 .muxIn_1(s_logisimBus7[31:0]),
                 .muxOut(s_logisimBus1[31:0]),
                 .sel(s_logisimBus6[31]));

   Multiplexer_bus_2 #(.nrOfBits(32))
      PLEXERS_2 (.enable(1'b1),
                 .muxIn_0(s_logisimBus8[31:0]),
                 .muxIn_1(s_logisimBus1[31:0]),
                 .muxOut(s_logisimBus6[63:32]),
                 .sel(s_logisimNet5));


endmodule
