/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
Onehot
**
**
**
*****************************************************************************/
module
Onehot(
Exec,
IDecode,
IFetch,
Instdone,
Mem,
WB,
clk,
rst
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
Instdone;
input
clk;
input
rst;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
Exec;
output
IDecode;
output
IFetch;
output
Mem;
output
WB;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
s_logisimNet0;
wire
s_logisimNet1;
wire
s_logisimNet10;
wire
s_logisimNet11;
wire
s_logisimNet2;
wire
s_logisimNet3;
wire
s_logisimNet4;
wire
s_logisimNet5;
wire
s_logisimNet6;
wire
s_logisimNet7;
wire
s_logisimNet8;
wire
s_logisimNet9;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimNet3
=
rst;
assign
s_logisimNet6
=
Instdone;
assign
s_logisimNet7
=
clk;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
Exec
=
s_logisimNet10;
assign
IDecode
=
s_logisimNet1;
assign
IFetch
=
s_logisimNet0;
assign
Mem
=
s_logisimNet11;
assign
WB
=
s_logisimNet5;
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimNet4
=
~s_logisimNet6;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
AND_GATE
#(.BubblesMask(2'b00))
GATES_1
(.input1(s_logisimNet4),
.input2(s_logisimNet10),
.result(s_logisimNet2));
AND_GATE
#(.BubblesMask(2'b00))
GATES_2
(.input1(s_logisimNet6),
.input2(s_logisimNet10),
.result(s_logisimNet9));
Multiplexer_2
PLEXERS_3
(.enable(1'b1),
.muxIn_0(s_logisimNet1),
.muxIn_1(s_logisimNet10),
.muxOut(s_logisimNet8),
.sel(s_logisimNet2));
D_FLIPFLOP
#(.invertClockEnable(0))
MEMORY_4
(.clock(s_logisimNet7),
.d(s_logisimNet5),
.preset(s_logisimNet3),
.q(s_logisimNet0),
.qBar(),
.reset(1'b0),
.tick(1'b1));
D_FLIPFLOP
#(.invertClockEnable(0))
MEMORY_5
(.clock(s_logisimNet7),
.d(s_logisimNet0),
.preset(1'b0),
.q(s_logisimNet1),
.qBar(),
.reset(s_logisimNet3),
.tick(1'b1));
D_FLIPFLOP
#(.invertClockEnable(0))
MEMORY_6
(.clock(s_logisimNet7),
.d(s_logisimNet8),
.preset(1'b0),
.q(s_logisimNet10),
.qBar(),
.reset(s_logisimNet3),
.tick(1'b1));
D_FLIPFLOP
#(.invertClockEnable(0))
MEMORY_7
(.clock(s_logisimNet7),
.d(s_logisimNet9),
.preset(1'b0),
.q(s_logisimNet11),
.qBar(),
.reset(s_logisimNet3),
.tick(1'b1));
D_FLIPFLOP
#(.invertClockEnable(0))
MEMORY_8
(.clock(s_logisimNet7),
.d(s_logisimNet11),
.preset(1'b0),
.q(s_logisimNet5),
.qBar(),
.reset(s_logisimNet3),
.tick(1'b1));
endmodule